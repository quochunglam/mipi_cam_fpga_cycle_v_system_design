// top.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module top (
		input  wire        clk_clk,                                                 //                                     clk.clk
		input  wire [2:0]  ddr3_status_external_connection_export,                  //         ddr3_status_external_connection.export
		input  wire [31:0] hip_ctrl_test_in,                                        //                                hip_ctrl.test_in
		input  wire        hip_ctrl_simu_mode_pipe,                                 //                                        .simu_mode_pipe
		input  wire        hip_pipe_sim_pipe_pclk_in,                               //                                hip_pipe.sim_pipe_pclk_in
		output wire [1:0]  hip_pipe_sim_pipe_rate,                                  //                                        .sim_pipe_rate
		output wire [4:0]  hip_pipe_sim_ltssmstate,                                 //                                        .sim_ltssmstate
		output wire [2:0]  hip_pipe_eidleinfersel0,                                 //                                        .eidleinfersel0
		output wire [2:0]  hip_pipe_eidleinfersel1,                                 //                                        .eidleinfersel1
		output wire [2:0]  hip_pipe_eidleinfersel2,                                 //                                        .eidleinfersel2
		output wire [2:0]  hip_pipe_eidleinfersel3,                                 //                                        .eidleinfersel3
		output wire [1:0]  hip_pipe_powerdown0,                                     //                                        .powerdown0
		output wire [1:0]  hip_pipe_powerdown1,                                     //                                        .powerdown1
		output wire [1:0]  hip_pipe_powerdown2,                                     //                                        .powerdown2
		output wire [1:0]  hip_pipe_powerdown3,                                     //                                        .powerdown3
		output wire        hip_pipe_rxpolarity0,                                    //                                        .rxpolarity0
		output wire        hip_pipe_rxpolarity1,                                    //                                        .rxpolarity1
		output wire        hip_pipe_rxpolarity2,                                    //                                        .rxpolarity2
		output wire        hip_pipe_rxpolarity3,                                    //                                        .rxpolarity3
		output wire        hip_pipe_txcompl0,                                       //                                        .txcompl0
		output wire        hip_pipe_txcompl1,                                       //                                        .txcompl1
		output wire        hip_pipe_txcompl2,                                       //                                        .txcompl2
		output wire        hip_pipe_txcompl3,                                       //                                        .txcompl3
		output wire [7:0]  hip_pipe_txdata0,                                        //                                        .txdata0
		output wire [7:0]  hip_pipe_txdata1,                                        //                                        .txdata1
		output wire [7:0]  hip_pipe_txdata2,                                        //                                        .txdata2
		output wire [7:0]  hip_pipe_txdata3,                                        //                                        .txdata3
		output wire        hip_pipe_txdatak0,                                       //                                        .txdatak0
		output wire        hip_pipe_txdatak1,                                       //                                        .txdatak1
		output wire        hip_pipe_txdatak2,                                       //                                        .txdatak2
		output wire        hip_pipe_txdatak3,                                       //                                        .txdatak3
		output wire        hip_pipe_txdetectrx0,                                    //                                        .txdetectrx0
		output wire        hip_pipe_txdetectrx1,                                    //                                        .txdetectrx1
		output wire        hip_pipe_txdetectrx2,                                    //                                        .txdetectrx2
		output wire        hip_pipe_txdetectrx3,                                    //                                        .txdetectrx3
		output wire        hip_pipe_txelecidle0,                                    //                                        .txelecidle0
		output wire        hip_pipe_txelecidle1,                                    //                                        .txelecidle1
		output wire        hip_pipe_txelecidle2,                                    //                                        .txelecidle2
		output wire        hip_pipe_txelecidle3,                                    //                                        .txelecidle3
		output wire        hip_pipe_txdeemph0,                                      //                                        .txdeemph0
		output wire        hip_pipe_txdeemph1,                                      //                                        .txdeemph1
		output wire        hip_pipe_txdeemph2,                                      //                                        .txdeemph2
		output wire        hip_pipe_txdeemph3,                                      //                                        .txdeemph3
		output wire [2:0]  hip_pipe_txmargin0,                                      //                                        .txmargin0
		output wire [2:0]  hip_pipe_txmargin1,                                      //                                        .txmargin1
		output wire [2:0]  hip_pipe_txmargin2,                                      //                                        .txmargin2
		output wire [2:0]  hip_pipe_txmargin3,                                      //                                        .txmargin3
		output wire        hip_pipe_txswing0,                                       //                                        .txswing0
		output wire        hip_pipe_txswing1,                                       //                                        .txswing1
		output wire        hip_pipe_txswing2,                                       //                                        .txswing2
		output wire        hip_pipe_txswing3,                                       //                                        .txswing3
		input  wire        hip_pipe_phystatus0,                                     //                                        .phystatus0
		input  wire        hip_pipe_phystatus1,                                     //                                        .phystatus1
		input  wire        hip_pipe_phystatus2,                                     //                                        .phystatus2
		input  wire        hip_pipe_phystatus3,                                     //                                        .phystatus3
		input  wire [7:0]  hip_pipe_rxdata0,                                        //                                        .rxdata0
		input  wire [7:0]  hip_pipe_rxdata1,                                        //                                        .rxdata1
		input  wire [7:0]  hip_pipe_rxdata2,                                        //                                        .rxdata2
		input  wire [7:0]  hip_pipe_rxdata3,                                        //                                        .rxdata3
		input  wire        hip_pipe_rxdatak0,                                       //                                        .rxdatak0
		input  wire        hip_pipe_rxdatak1,                                       //                                        .rxdatak1
		input  wire        hip_pipe_rxdatak2,                                       //                                        .rxdatak2
		input  wire        hip_pipe_rxdatak3,                                       //                                        .rxdatak3
		input  wire        hip_pipe_rxelecidle0,                                    //                                        .rxelecidle0
		input  wire        hip_pipe_rxelecidle1,                                    //                                        .rxelecidle1
		input  wire        hip_pipe_rxelecidle2,                                    //                                        .rxelecidle2
		input  wire        hip_pipe_rxelecidle3,                                    //                                        .rxelecidle3
		input  wire [2:0]  hip_pipe_rxstatus0,                                      //                                        .rxstatus0
		input  wire [2:0]  hip_pipe_rxstatus1,                                      //                                        .rxstatus1
		input  wire [2:0]  hip_pipe_rxstatus2,                                      //                                        .rxstatus2
		input  wire [2:0]  hip_pipe_rxstatus3,                                      //                                        .rxstatus3
		input  wire        hip_pipe_rxvalid0,                                       //                                        .rxvalid0
		input  wire        hip_pipe_rxvalid1,                                       //                                        .rxvalid1
		input  wire        hip_pipe_rxvalid2,                                       //                                        .rxvalid2
		input  wire        hip_pipe_rxvalid3,                                       //                                        .rxvalid3
		input  wire        hip_serial_rx_in0,                                       //                              hip_serial.rx_in0
		input  wire        hip_serial_rx_in1,                                       //                                        .rx_in1
		input  wire        hip_serial_rx_in2,                                       //                                        .rx_in2
		input  wire        hip_serial_rx_in3,                                       //                                        .rx_in3
		output wire        hip_serial_tx_out0,                                      //                                        .tx_out0
		output wire        hip_serial_tx_out1,                                      //                                        .tx_out1
		output wire        hip_serial_tx_out2,                                      //                                        .tx_out2
		output wire        hip_serial_tx_out3,                                      //                                        .tx_out3
		inout  wire        i2c_opencores_camera_export_scl_pad_io,                  //             i2c_opencores_camera_export.scl_pad_io
		inout  wire        i2c_opencores_camera_export_sda_pad_io,                  //                                        .sda_pad_io
		inout  wire        i2c_opencores_mipi_export_scl_pad_io,                    //               i2c_opencores_mipi_export.scl_pad_io
		inout  wire        i2c_opencores_mipi_export_sda_pad_io,                    //                                        .sda_pad_io
		input  wire        mem_if_ddr3_emif_0_pll_ref_clk_clk,                      //          mem_if_ddr3_emif_0_pll_ref_clk.clk
		output wire        mem_if_ddr3_emif_0_status_local_init_done,               //               mem_if_ddr3_emif_0_status.local_init_done
		output wire        mem_if_ddr3_emif_0_status_local_cal_success,             //                                        .local_cal_success
		output wire        mem_if_ddr3_emif_0_status_local_cal_fail,                //                                        .local_cal_fail
		output wire [14:0] memory_mem_a,                                            //                                  memory.mem_a
		output wire [2:0]  memory_mem_ba,                                           //                                        .mem_ba
		output wire [0:0]  memory_mem_ck,                                           //                                        .mem_ck
		output wire [0:0]  memory_mem_ck_n,                                         //                                        .mem_ck_n
		output wire [0:0]  memory_mem_cke,                                          //                                        .mem_cke
		output wire [0:0]  memory_mem_cs_n,                                         //                                        .mem_cs_n
		output wire [3:0]  memory_mem_dm,                                           //                                        .mem_dm
		output wire [0:0]  memory_mem_ras_n,                                        //                                        .mem_ras_n
		output wire [0:0]  memory_mem_cas_n,                                        //                                        .mem_cas_n
		output wire [0:0]  memory_mem_we_n,                                         //                                        .mem_we_n
		output wire        memory_mem_reset_n,                                      //                                        .mem_reset_n
		inout  wire [31:0] memory_mem_dq,                                           //                                        .mem_dq
		inout  wire [3:0]  memory_mem_dqs,                                          //                                        .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,                                        //                                        .mem_dqs_n
		output wire [0:0]  memory_mem_odt,                                          //                                        .mem_odt
		output wire        mipi_pwdn_n_external_connection_export,                  //         mipi_pwdn_n_external_connection.export
		output wire        mipi_reset_n_external_connection_export,                 //        mipi_reset_n_external_connection.export
		input  wire        oct_rzqin,                                               //                                     oct.rzqin
		output wire        pcie_256_hip_avmm_0_reconfig_clk_locked_fixedclk_locked, // pcie_256_hip_avmm_0_reconfig_clk_locked.fixedclk_locked
		input  wire        pcie_rstn_npor,                                          //                               pcie_rstn.npor
		input  wire        pcie_rstn_pin_perst,                                     //                                        .pin_perst
		input  wire [3:0]  pio_button_external_connection_export,                   //          pio_button_external_connection.export
		output wire [3:0]  pio_led_external_connection_export,                      //             pio_led_external_connection.export
		output wire        pll_0_outclk1_100mhz_clk,                                //                    pll_0_outclk1_100mhz.clk
		output wire        pll_0_outclk2_20mhz_clk,                                 //                     pll_0_outclk2_20mhz.clk
		input  wire        refclk_clk,                                              //                                  refclk.clk
		input  wire        reset_reset_n,                                           //                                   reset.reset_n
		output wire [12:0] sdram_vfb_wire_addr,                                     //                          sdram_vfb_wire.addr
		output wire [1:0]  sdram_vfb_wire_ba,                                       //                                        .ba
		output wire        sdram_vfb_wire_cas_n,                                    //                                        .cas_n
		output wire        sdram_vfb_wire_cke,                                      //                                        .cke
		output wire        sdram_vfb_wire_cs_n,                                     //                                        .cs_n
		inout  wire [15:0] sdram_vfb_wire_dq,                                       //                                        .dq
		output wire [1:0]  sdram_vfb_wire_dqm,                                      //                                        .dqm
		output wire        sdram_vfb_wire_ras_n,                                    //                                        .ras_n
		output wire        sdram_vfb_wire_we_n,                                     //                                        .we_n
		inout  wire        terasic_auto_focus_0_conduit_vcm_i2c_sda,                //            terasic_auto_focus_0_conduit.vcm_i2c_sda
		input  wire        terasic_auto_focus_0_conduit_clk50,                      //                                        .clk50
		inout  wire        terasic_auto_focus_0_conduit_vcm_i2c_scl,                //                                        .vcm_i2c_scl
		input  wire [11:0] terasic_camera_0_conduit_end_cam_d,                      //            terasic_camera_0_conduit_end.cam_d
		input  wire        terasic_camera_0_conduit_end_cam_fval,                   //                                        .cam_fval
		input  wire        terasic_camera_0_conduit_end_cam_lval,                   //                                        .cam_lval
		input  wire        terasic_camera_0_conduit_end_cam_pix                     //                                        .cam_pix
	);

	wire          alt_vip_cl_vfb_0_dout_valid;                                       // alt_vip_cl_vfb_0:dout_valid -> TERASIC_AUTO_FOCUS_0:sink_valid
	wire   [23:0] alt_vip_cl_vfb_0_dout_data;                                        // alt_vip_cl_vfb_0:dout_data -> TERASIC_AUTO_FOCUS_0:sink_data
	wire          alt_vip_cl_vfb_0_dout_ready;                                       // TERASIC_AUTO_FOCUS_0:sink_ready -> alt_vip_cl_vfb_0:dout_ready
	wire          alt_vip_cl_vfb_0_dout_startofpacket;                               // alt_vip_cl_vfb_0:dout_startofpacket -> TERASIC_AUTO_FOCUS_0:sink_sop
	wire          alt_vip_cl_vfb_0_dout_endofpacket;                                 // alt_vip_cl_vfb_0:dout_endofpacket -> TERASIC_AUTO_FOCUS_0:sink_eop
	wire          pcie_256_dma_coreclkout_clk;                                       // pcie_256_dma:coreclkout -> [csr_regmap:clk2, mm_interconnect_0:pcie_256_dma_coreclkout_clk, mm_interconnect_2:pcie_256_dma_coreclkout_clk, mm_interconnect_4:pcie_256_dma_coreclkout_clk, mm_interconnect_5:pcie_256_dma_coreclkout_clk, ocm_256k_dma:clk2, pcie_reconfig_driver_0:pld_clk, pcie_reconfig_driver_0:reconfig_xcvr_clk, rst_controller_002:clk]
	wire          pll_0_outclk0_clk;                                                 // pll_0:outclk_0 -> [TERASIC_AUTO_FOCUS_0:clk, TERASIC_CAMERA_0:clk, alt_vip_cl_vfb_0:main_clock, avalon_st_adapter:in_clk_0_clk, avalon_st_adapter_001:in_clk_0_clk, csr_regmap:clk, ddr3_status:clk, fifo_0:wrclock, i2c_opencores_camera:wb_clk_i, i2c_opencores_mipi:wb_clk_i, irq_mapper:clk, jtag_uart_0:clk, mem_if_ddr3_emif_0:mp_cmd_clk_0_clk, mem_if_ddr3_emif_0:mp_rfifo_clk_0_clk, mem_if_ddr3_emif_0:mp_rfifo_clk_1_clk, mem_if_ddr3_emif_0:mp_wfifo_clk_0_clk, mem_if_ddr3_emif_0:mp_wfifo_clk_1_clk, mipi_pwdn_n:clk, mipi_reset_n:clk, mm_interconnect_1:pll_0_outclk0_clk, mm_interconnect_3:pll_0_outclk0_clk, nios2_gen2_0:clk, nios_ram:clk, ocm_256k_dma:clk, pio_button:clk, pio_led:clk, rst_controller:clk, sdram_vfb:clk, sysid_qsys_0:clock, timer_0:clk]
	wire    [1:0] pcie_256_dma_hip_currentspeed_currentspeed;                        // pcie_256_dma:currentspeed -> pcie_reconfig_driver_0:currentspeed
	wire  [229:0] pcie_256_dma_reconfig_from_xcvr_reconfig_from_xcvr;                // pcie_256_dma:reconfig_from_xcvr -> alt_xcvr_reconfig_0:reconfig_from_xcvr
	wire  [349:0] alt_xcvr_reconfig_0_reconfig_to_xcvr_reconfig_to_xcvr;             // alt_xcvr_reconfig_0:reconfig_to_xcvr -> pcie_256_dma:reconfig_to_xcvr
	wire          pcie_256_dma_rxm_bar2_waitrequest;                                 // mm_interconnect_0:pcie_256_dma_Rxm_BAR2_waitrequest -> pcie_256_dma:RxmWaitRequest_2_i
	wire   [31:0] pcie_256_dma_rxm_bar2_readdata;                                    // mm_interconnect_0:pcie_256_dma_Rxm_BAR2_readdata -> pcie_256_dma:RxmReadData_2_i
	wire   [63:0] pcie_256_dma_rxm_bar2_address;                                     // pcie_256_dma:RxmAddress_2_o -> mm_interconnect_0:pcie_256_dma_Rxm_BAR2_address
	wire          pcie_256_dma_rxm_bar2_read;                                        // pcie_256_dma:RxmRead_2_o -> mm_interconnect_0:pcie_256_dma_Rxm_BAR2_read
	wire    [3:0] pcie_256_dma_rxm_bar2_byteenable;                                  // pcie_256_dma:RxmByteEnable_2_o -> mm_interconnect_0:pcie_256_dma_Rxm_BAR2_byteenable
	wire          pcie_256_dma_rxm_bar2_readdatavalid;                               // mm_interconnect_0:pcie_256_dma_Rxm_BAR2_readdatavalid -> pcie_256_dma:RxmReadDataValid_2_i
	wire          pcie_256_dma_rxm_bar2_write;                                       // pcie_256_dma:RxmWrite_2_o -> mm_interconnect_0:pcie_256_dma_Rxm_BAR2_write
	wire   [31:0] pcie_256_dma_rxm_bar2_writedata;                                   // pcie_256_dma:RxmWriteData_2_o -> mm_interconnect_0:pcie_256_dma_Rxm_BAR2_writedata
	wire          mm_interconnect_0_csr_regmap_s2_chipselect;                        // mm_interconnect_0:csr_regmap_s2_chipselect -> csr_regmap:chipselect2
	wire   [31:0] mm_interconnect_0_csr_regmap_s2_readdata;                          // csr_regmap:readdata2 -> mm_interconnect_0:csr_regmap_s2_readdata
	wire    [2:0] mm_interconnect_0_csr_regmap_s2_address;                           // mm_interconnect_0:csr_regmap_s2_address -> csr_regmap:address2
	wire    [3:0] mm_interconnect_0_csr_regmap_s2_byteenable;                        // mm_interconnect_0:csr_regmap_s2_byteenable -> csr_regmap:byteenable2
	wire          mm_interconnect_0_csr_regmap_s2_write;                             // mm_interconnect_0:csr_regmap_s2_write -> csr_regmap:write2
	wire   [31:0] mm_interconnect_0_csr_regmap_s2_writedata;                         // mm_interconnect_0:csr_regmap_s2_writedata -> csr_regmap:writedata2
	wire          mm_interconnect_0_csr_regmap_s2_clken;                             // mm_interconnect_0:csr_regmap_s2_clken -> csr_regmap:clken2
	wire   [31:0] nios2_gen2_0_data_master_readdata;                                 // mm_interconnect_1:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire          nios2_gen2_0_data_master_waitrequest;                              // mm_interconnect_1:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire          nios2_gen2_0_data_master_debugaccess;                              // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_1:nios2_gen2_0_data_master_debugaccess
	wire   [30:0] nios2_gen2_0_data_master_address;                                  // nios2_gen2_0:d_address -> mm_interconnect_1:nios2_gen2_0_data_master_address
	wire    [3:0] nios2_gen2_0_data_master_byteenable;                               // nios2_gen2_0:d_byteenable -> mm_interconnect_1:nios2_gen2_0_data_master_byteenable
	wire          nios2_gen2_0_data_master_read;                                     // nios2_gen2_0:d_read -> mm_interconnect_1:nios2_gen2_0_data_master_read
	wire          nios2_gen2_0_data_master_readdatavalid;                            // mm_interconnect_1:nios2_gen2_0_data_master_readdatavalid -> nios2_gen2_0:d_readdatavalid
	wire          nios2_gen2_0_data_master_write;                                    // nios2_gen2_0:d_write -> mm_interconnect_1:nios2_gen2_0_data_master_write
	wire   [31:0] nios2_gen2_0_data_master_writedata;                                // nios2_gen2_0:d_writedata -> mm_interconnect_1:nios2_gen2_0_data_master_writedata
	wire   [31:0] nios2_gen2_0_instruction_master_readdata;                          // mm_interconnect_1:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire          nios2_gen2_0_instruction_master_waitrequest;                       // mm_interconnect_1:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire   [30:0] nios2_gen2_0_instruction_master_address;                           // nios2_gen2_0:i_address -> mm_interconnect_1:nios2_gen2_0_instruction_master_address
	wire          nios2_gen2_0_instruction_master_read;                              // nios2_gen2_0:i_read -> mm_interconnect_1:nios2_gen2_0_instruction_master_read
	wire          nios2_gen2_0_instruction_master_readdatavalid;                     // mm_interconnect_1:nios2_gen2_0_instruction_master_readdatavalid -> nios2_gen2_0:i_readdatavalid
	wire          mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_chipselect;        // mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire   [31:0] mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_readdata;          // jtag_uart_0:av_readdata -> mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_readdata
	wire          mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_waitrequest;       // jtag_uart_0:av_waitrequest -> mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire    [0:0] mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_address;           // mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire          mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read;              // mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire          mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write;             // mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire   [31:0] mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_writedata;         // mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire          mm_interconnect_1_i2c_opencores_camera_avalon_slave_0_chipselect;  // mm_interconnect_1:i2c_opencores_camera_avalon_slave_0_chipselect -> i2c_opencores_camera:wb_stb_i
	wire    [7:0] mm_interconnect_1_i2c_opencores_camera_avalon_slave_0_readdata;    // i2c_opencores_camera:wb_dat_o -> mm_interconnect_1:i2c_opencores_camera_avalon_slave_0_readdata
	wire          mm_interconnect_1_i2c_opencores_camera_avalon_slave_0_waitrequest; // i2c_opencores_camera:wb_ack_o -> mm_interconnect_1:i2c_opencores_camera_avalon_slave_0_waitrequest
	wire    [2:0] mm_interconnect_1_i2c_opencores_camera_avalon_slave_0_address;     // mm_interconnect_1:i2c_opencores_camera_avalon_slave_0_address -> i2c_opencores_camera:wb_adr_i
	wire          mm_interconnect_1_i2c_opencores_camera_avalon_slave_0_write;       // mm_interconnect_1:i2c_opencores_camera_avalon_slave_0_write -> i2c_opencores_camera:wb_we_i
	wire    [7:0] mm_interconnect_1_i2c_opencores_camera_avalon_slave_0_writedata;   // mm_interconnect_1:i2c_opencores_camera_avalon_slave_0_writedata -> i2c_opencores_camera:wb_dat_i
	wire          mm_interconnect_1_i2c_opencores_mipi_avalon_slave_0_chipselect;    // mm_interconnect_1:i2c_opencores_mipi_avalon_slave_0_chipselect -> i2c_opencores_mipi:wb_stb_i
	wire    [7:0] mm_interconnect_1_i2c_opencores_mipi_avalon_slave_0_readdata;      // i2c_opencores_mipi:wb_dat_o -> mm_interconnect_1:i2c_opencores_mipi_avalon_slave_0_readdata
	wire          mm_interconnect_1_i2c_opencores_mipi_avalon_slave_0_waitrequest;   // i2c_opencores_mipi:wb_ack_o -> mm_interconnect_1:i2c_opencores_mipi_avalon_slave_0_waitrequest
	wire    [2:0] mm_interconnect_1_i2c_opencores_mipi_avalon_slave_0_address;       // mm_interconnect_1:i2c_opencores_mipi_avalon_slave_0_address -> i2c_opencores_mipi:wb_adr_i
	wire          mm_interconnect_1_i2c_opencores_mipi_avalon_slave_0_write;         // mm_interconnect_1:i2c_opencores_mipi_avalon_slave_0_write -> i2c_opencores_mipi:wb_we_i
	wire    [7:0] mm_interconnect_1_i2c_opencores_mipi_avalon_slave_0_writedata;     // mm_interconnect_1:i2c_opencores_mipi_avalon_slave_0_writedata -> i2c_opencores_mipi:wb_dat_i
	wire          mm_interconnect_1_mem_if_ddr3_emif_0_avl_0_beginbursttransfer;     // mm_interconnect_1:mem_if_ddr3_emif_0_avl_0_beginbursttransfer -> mem_if_ddr3_emif_0:avl_burstbegin_0
	wire  [127:0] mm_interconnect_1_mem_if_ddr3_emif_0_avl_0_readdata;               // mem_if_ddr3_emif_0:avl_rdata_0 -> mm_interconnect_1:mem_if_ddr3_emif_0_avl_0_readdata
	wire          mm_interconnect_1_mem_if_ddr3_emif_0_avl_0_waitrequest;            // mem_if_ddr3_emif_0:avl_ready_0 -> mm_interconnect_1:mem_if_ddr3_emif_0_avl_0_waitrequest
	wire   [25:0] mm_interconnect_1_mem_if_ddr3_emif_0_avl_0_address;                // mm_interconnect_1:mem_if_ddr3_emif_0_avl_0_address -> mem_if_ddr3_emif_0:avl_addr_0
	wire          mm_interconnect_1_mem_if_ddr3_emif_0_avl_0_read;                   // mm_interconnect_1:mem_if_ddr3_emif_0_avl_0_read -> mem_if_ddr3_emif_0:avl_read_req_0
	wire   [15:0] mm_interconnect_1_mem_if_ddr3_emif_0_avl_0_byteenable;             // mm_interconnect_1:mem_if_ddr3_emif_0_avl_0_byteenable -> mem_if_ddr3_emif_0:avl_be_0
	wire          mm_interconnect_1_mem_if_ddr3_emif_0_avl_0_readdatavalid;          // mem_if_ddr3_emif_0:avl_rdata_valid_0 -> mm_interconnect_1:mem_if_ddr3_emif_0_avl_0_readdatavalid
	wire          mm_interconnect_1_mem_if_ddr3_emif_0_avl_0_write;                  // mm_interconnect_1:mem_if_ddr3_emif_0_avl_0_write -> mem_if_ddr3_emif_0:avl_write_req_0
	wire  [127:0] mm_interconnect_1_mem_if_ddr3_emif_0_avl_0_writedata;              // mm_interconnect_1:mem_if_ddr3_emif_0_avl_0_writedata -> mem_if_ddr3_emif_0:avl_wdata_0
	wire    [5:0] mm_interconnect_1_mem_if_ddr3_emif_0_avl_0_burstcount;             // mm_interconnect_1:mem_if_ddr3_emif_0_avl_0_burstcount -> mem_if_ddr3_emif_0:avl_size_0
	wire   [31:0] mm_interconnect_1_sysid_qsys_0_control_slave_readdata;             // sysid_qsys_0:readdata -> mm_interconnect_1:sysid_qsys_0_control_slave_readdata
	wire    [0:0] mm_interconnect_1_sysid_qsys_0_control_slave_address;              // mm_interconnect_1:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire   [31:0] mm_interconnect_1_nios2_gen2_0_debug_mem_slave_readdata;           // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_1:nios2_gen2_0_debug_mem_slave_readdata
	wire          mm_interconnect_1_nios2_gen2_0_debug_mem_slave_waitrequest;        // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_1:nios2_gen2_0_debug_mem_slave_waitrequest
	wire          mm_interconnect_1_nios2_gen2_0_debug_mem_slave_debugaccess;        // mm_interconnect_1:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire    [8:0] mm_interconnect_1_nios2_gen2_0_debug_mem_slave_address;            // mm_interconnect_1:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire          mm_interconnect_1_nios2_gen2_0_debug_mem_slave_read;               // mm_interconnect_1:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire    [3:0] mm_interconnect_1_nios2_gen2_0_debug_mem_slave_byteenable;         // mm_interconnect_1:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire          mm_interconnect_1_nios2_gen2_0_debug_mem_slave_write;              // mm_interconnect_1:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire   [31:0] mm_interconnect_1_nios2_gen2_0_debug_mem_slave_writedata;          // mm_interconnect_1:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire   [31:0] mm_interconnect_1_fifo_0_in_csr_readdata;                          // fifo_0:wrclk_control_slave_readdata -> mm_interconnect_1:fifo_0_in_csr_readdata
	wire    [2:0] mm_interconnect_1_fifo_0_in_csr_address;                           // mm_interconnect_1:fifo_0_in_csr_address -> fifo_0:wrclk_control_slave_address
	wire          mm_interconnect_1_fifo_0_in_csr_read;                              // mm_interconnect_1:fifo_0_in_csr_read -> fifo_0:wrclk_control_slave_read
	wire          mm_interconnect_1_fifo_0_in_csr_write;                             // mm_interconnect_1:fifo_0_in_csr_write -> fifo_0:wrclk_control_slave_write
	wire   [31:0] mm_interconnect_1_fifo_0_in_csr_writedata;                         // mm_interconnect_1:fifo_0_in_csr_writedata -> fifo_0:wrclk_control_slave_writedata
	wire          mm_interconnect_1_terasic_auto_focus_0_mm_ctrl_chipselect;         // mm_interconnect_1:TERASIC_AUTO_FOCUS_0_mm_ctrl_chipselect -> TERASIC_AUTO_FOCUS_0:s_chipselect
	wire   [31:0] mm_interconnect_1_terasic_auto_focus_0_mm_ctrl_readdata;           // TERASIC_AUTO_FOCUS_0:s_readdata -> mm_interconnect_1:TERASIC_AUTO_FOCUS_0_mm_ctrl_readdata
	wire    [2:0] mm_interconnect_1_terasic_auto_focus_0_mm_ctrl_address;            // mm_interconnect_1:TERASIC_AUTO_FOCUS_0_mm_ctrl_address -> TERASIC_AUTO_FOCUS_0:s_address
	wire          mm_interconnect_1_terasic_auto_focus_0_mm_ctrl_read;               // mm_interconnect_1:TERASIC_AUTO_FOCUS_0_mm_ctrl_read -> TERASIC_AUTO_FOCUS_0:s_read
	wire          mm_interconnect_1_terasic_auto_focus_0_mm_ctrl_write;              // mm_interconnect_1:TERASIC_AUTO_FOCUS_0_mm_ctrl_write -> TERASIC_AUTO_FOCUS_0:s_write
	wire   [31:0] mm_interconnect_1_terasic_auto_focus_0_mm_ctrl_writedata;          // mm_interconnect_1:TERASIC_AUTO_FOCUS_0_mm_ctrl_writedata -> TERASIC_AUTO_FOCUS_0:s_writedata
	wire   [31:0] mm_interconnect_1_fifo_0_out_readdata;                             // fifo_0:avalonmm_read_slave_readdata -> mm_interconnect_1:fifo_0_out_readdata
	wire          mm_interconnect_1_fifo_0_out_waitrequest;                          // fifo_0:avalonmm_read_slave_waitrequest -> mm_interconnect_1:fifo_0_out_waitrequest
	wire    [0:0] mm_interconnect_1_fifo_0_out_address;                              // mm_interconnect_1:fifo_0_out_address -> fifo_0:avalonmm_read_slave_address
	wire          mm_interconnect_1_fifo_0_out_read;                                 // mm_interconnect_1:fifo_0_out_read -> fifo_0:avalonmm_read_slave_read
	wire          mm_interconnect_1_nios_ram_s1_chipselect;                          // mm_interconnect_1:nios_ram_s1_chipselect -> nios_ram:chipselect
	wire   [31:0] mm_interconnect_1_nios_ram_s1_readdata;                            // nios_ram:readdata -> mm_interconnect_1:nios_ram_s1_readdata
	wire   [14:0] mm_interconnect_1_nios_ram_s1_address;                             // mm_interconnect_1:nios_ram_s1_address -> nios_ram:address
	wire    [3:0] mm_interconnect_1_nios_ram_s1_byteenable;                          // mm_interconnect_1:nios_ram_s1_byteenable -> nios_ram:byteenable
	wire          mm_interconnect_1_nios_ram_s1_write;                               // mm_interconnect_1:nios_ram_s1_write -> nios_ram:write
	wire   [31:0] mm_interconnect_1_nios_ram_s1_writedata;                           // mm_interconnect_1:nios_ram_s1_writedata -> nios_ram:writedata
	wire          mm_interconnect_1_nios_ram_s1_clken;                               // mm_interconnect_1:nios_ram_s1_clken -> nios_ram:clken
	wire          mm_interconnect_1_pio_led_s1_chipselect;                           // mm_interconnect_1:pio_led_s1_chipselect -> pio_led:chipselect
	wire   [31:0] mm_interconnect_1_pio_led_s1_readdata;                             // pio_led:readdata -> mm_interconnect_1:pio_led_s1_readdata
	wire    [1:0] mm_interconnect_1_pio_led_s1_address;                              // mm_interconnect_1:pio_led_s1_address -> pio_led:address
	wire          mm_interconnect_1_pio_led_s1_write;                                // mm_interconnect_1:pio_led_s1_write -> pio_led:write_n
	wire   [31:0] mm_interconnect_1_pio_led_s1_writedata;                            // mm_interconnect_1:pio_led_s1_writedata -> pio_led:writedata
	wire          mm_interconnect_1_pio_button_s1_chipselect;                        // mm_interconnect_1:pio_button_s1_chipselect -> pio_button:chipselect
	wire   [31:0] mm_interconnect_1_pio_button_s1_readdata;                          // pio_button:readdata -> mm_interconnect_1:pio_button_s1_readdata
	wire    [1:0] mm_interconnect_1_pio_button_s1_address;                           // mm_interconnect_1:pio_button_s1_address -> pio_button:address
	wire          mm_interconnect_1_pio_button_s1_write;                             // mm_interconnect_1:pio_button_s1_write -> pio_button:write_n
	wire   [31:0] mm_interconnect_1_pio_button_s1_writedata;                         // mm_interconnect_1:pio_button_s1_writedata -> pio_button:writedata
	wire          mm_interconnect_1_mipi_reset_n_s1_chipselect;                      // mm_interconnect_1:mipi_reset_n_s1_chipselect -> mipi_reset_n:chipselect
	wire   [31:0] mm_interconnect_1_mipi_reset_n_s1_readdata;                        // mipi_reset_n:readdata -> mm_interconnect_1:mipi_reset_n_s1_readdata
	wire    [1:0] mm_interconnect_1_mipi_reset_n_s1_address;                         // mm_interconnect_1:mipi_reset_n_s1_address -> mipi_reset_n:address
	wire          mm_interconnect_1_mipi_reset_n_s1_write;                           // mm_interconnect_1:mipi_reset_n_s1_write -> mipi_reset_n:write_n
	wire   [31:0] mm_interconnect_1_mipi_reset_n_s1_writedata;                       // mm_interconnect_1:mipi_reset_n_s1_writedata -> mipi_reset_n:writedata
	wire          mm_interconnect_1_mipi_pwdn_n_s1_chipselect;                       // mm_interconnect_1:mipi_pwdn_n_s1_chipselect -> mipi_pwdn_n:chipselect
	wire   [31:0] mm_interconnect_1_mipi_pwdn_n_s1_readdata;                         // mipi_pwdn_n:readdata -> mm_interconnect_1:mipi_pwdn_n_s1_readdata
	wire    [1:0] mm_interconnect_1_mipi_pwdn_n_s1_address;                          // mm_interconnect_1:mipi_pwdn_n_s1_address -> mipi_pwdn_n:address
	wire          mm_interconnect_1_mipi_pwdn_n_s1_write;                            // mm_interconnect_1:mipi_pwdn_n_s1_write -> mipi_pwdn_n:write_n
	wire   [31:0] mm_interconnect_1_mipi_pwdn_n_s1_writedata;                        // mm_interconnect_1:mipi_pwdn_n_s1_writedata -> mipi_pwdn_n:writedata
	wire          mm_interconnect_1_timer_0_s1_chipselect;                           // mm_interconnect_1:timer_0_s1_chipselect -> timer_0:chipselect
	wire   [15:0] mm_interconnect_1_timer_0_s1_readdata;                             // timer_0:readdata -> mm_interconnect_1:timer_0_s1_readdata
	wire    [2:0] mm_interconnect_1_timer_0_s1_address;                              // mm_interconnect_1:timer_0_s1_address -> timer_0:address
	wire          mm_interconnect_1_timer_0_s1_write;                                // mm_interconnect_1:timer_0_s1_write -> timer_0:write_n
	wire   [15:0] mm_interconnect_1_timer_0_s1_writedata;                            // mm_interconnect_1:timer_0_s1_writedata -> timer_0:writedata
	wire          mm_interconnect_1_ocm_256k_dma_s1_chipselect;                      // mm_interconnect_1:ocm_256k_dma_s1_chipselect -> ocm_256k_dma:chipselect
	wire   [31:0] mm_interconnect_1_ocm_256k_dma_s1_readdata;                        // ocm_256k_dma:readdata -> mm_interconnect_1:ocm_256k_dma_s1_readdata
	wire   [15:0] mm_interconnect_1_ocm_256k_dma_s1_address;                         // mm_interconnect_1:ocm_256k_dma_s1_address -> ocm_256k_dma:address
	wire    [3:0] mm_interconnect_1_ocm_256k_dma_s1_byteenable;                      // mm_interconnect_1:ocm_256k_dma_s1_byteenable -> ocm_256k_dma:byteenable
	wire          mm_interconnect_1_ocm_256k_dma_s1_write;                           // mm_interconnect_1:ocm_256k_dma_s1_write -> ocm_256k_dma:write
	wire   [31:0] mm_interconnect_1_ocm_256k_dma_s1_writedata;                       // mm_interconnect_1:ocm_256k_dma_s1_writedata -> ocm_256k_dma:writedata
	wire          mm_interconnect_1_ocm_256k_dma_s1_clken;                           // mm_interconnect_1:ocm_256k_dma_s1_clken -> ocm_256k_dma:clken
	wire          mm_interconnect_1_csr_regmap_s1_chipselect;                        // mm_interconnect_1:csr_regmap_s1_chipselect -> csr_regmap:chipselect
	wire   [31:0] mm_interconnect_1_csr_regmap_s1_readdata;                          // csr_regmap:readdata -> mm_interconnect_1:csr_regmap_s1_readdata
	wire    [2:0] mm_interconnect_1_csr_regmap_s1_address;                           // mm_interconnect_1:csr_regmap_s1_address -> csr_regmap:address
	wire    [3:0] mm_interconnect_1_csr_regmap_s1_byteenable;                        // mm_interconnect_1:csr_regmap_s1_byteenable -> csr_regmap:byteenable
	wire          mm_interconnect_1_csr_regmap_s1_write;                             // mm_interconnect_1:csr_regmap_s1_write -> csr_regmap:write
	wire   [31:0] mm_interconnect_1_csr_regmap_s1_writedata;                         // mm_interconnect_1:csr_regmap_s1_writedata -> csr_regmap:writedata
	wire          mm_interconnect_1_csr_regmap_s1_clken;                             // mm_interconnect_1:csr_regmap_s1_clken -> csr_regmap:clken
	wire   [31:0] mm_interconnect_1_ddr3_status_s1_readdata;                         // ddr3_status:readdata -> mm_interconnect_1:ddr3_status_s1_readdata
	wire    [1:0] mm_interconnect_1_ddr3_status_s1_address;                          // mm_interconnect_1:ddr3_status_s1_address -> ddr3_status:address
	wire          pcie_256_dma_dma_rd_master_waitrequest;                            // mm_interconnect_2:pcie_256_dma_dma_rd_master_waitrequest -> pcie_256_dma:RdDmaWaitRequest_i
	wire   [63:0] pcie_256_dma_dma_rd_master_address;                                // pcie_256_dma:RdDmaAddress_o -> mm_interconnect_2:pcie_256_dma_dma_rd_master_address
	wire   [15:0] pcie_256_dma_dma_rd_master_byteenable;                             // pcie_256_dma:RdDmaWriteEnable_o -> mm_interconnect_2:pcie_256_dma_dma_rd_master_byteenable
	wire          pcie_256_dma_dma_rd_master_write;                                  // pcie_256_dma:RdDmaWrite_o -> mm_interconnect_2:pcie_256_dma_dma_rd_master_write
	wire  [127:0] pcie_256_dma_dma_rd_master_writedata;                              // pcie_256_dma:RdDmaWriteData_o -> mm_interconnect_2:pcie_256_dma_dma_rd_master_writedata
	wire    [5:0] pcie_256_dma_dma_rd_master_burstcount;                             // pcie_256_dma:RdDmaBurstCount_o -> mm_interconnect_2:pcie_256_dma_dma_rd_master_burstcount
	wire          pcie_256_dma_dma_wr_master_waitrequest;                            // mm_interconnect_2:pcie_256_dma_dma_wr_master_waitrequest -> pcie_256_dma:WrDmaWaitRequest_i
	wire  [127:0] pcie_256_dma_dma_wr_master_readdata;                               // mm_interconnect_2:pcie_256_dma_dma_wr_master_readdata -> pcie_256_dma:WrDmaReadData_i
	wire   [63:0] pcie_256_dma_dma_wr_master_address;                                // pcie_256_dma:WrDmaAddress_o -> mm_interconnect_2:pcie_256_dma_dma_wr_master_address
	wire          pcie_256_dma_dma_wr_master_read;                                   // pcie_256_dma:WrDmaRead_o -> mm_interconnect_2:pcie_256_dma_dma_wr_master_read
	wire          pcie_256_dma_dma_wr_master_readdatavalid;                          // mm_interconnect_2:pcie_256_dma_dma_wr_master_readdatavalid -> pcie_256_dma:WrDmaReadDataValid_i
	wire    [5:0] pcie_256_dma_dma_wr_master_burstcount;                             // pcie_256_dma:WrDmaBurstCount_o -> mm_interconnect_2:pcie_256_dma_dma_wr_master_burstcount
	wire          mm_interconnect_2_pcie_256_dma_rd_dts_slave_chipselect;            // mm_interconnect_2:pcie_256_dma_rd_dts_slave_chipselect -> pcie_256_dma:RdDTSChipSelect_i
	wire          mm_interconnect_2_pcie_256_dma_rd_dts_slave_waitrequest;           // pcie_256_dma:RdDTSWaitRequest_o -> mm_interconnect_2:pcie_256_dma_rd_dts_slave_waitrequest
	wire    [7:0] mm_interconnect_2_pcie_256_dma_rd_dts_slave_address;               // mm_interconnect_2:pcie_256_dma_rd_dts_slave_address -> pcie_256_dma:RdDTSAddress_i
	wire          mm_interconnect_2_pcie_256_dma_rd_dts_slave_write;                 // mm_interconnect_2:pcie_256_dma_rd_dts_slave_write -> pcie_256_dma:RdDTSWrite_i
	wire  [255:0] mm_interconnect_2_pcie_256_dma_rd_dts_slave_writedata;             // mm_interconnect_2:pcie_256_dma_rd_dts_slave_writedata -> pcie_256_dma:RdDTSWriteData_i
	wire    [4:0] mm_interconnect_2_pcie_256_dma_rd_dts_slave_burstcount;            // mm_interconnect_2:pcie_256_dma_rd_dts_slave_burstcount -> pcie_256_dma:RdDTSBurstCount_i
	wire          mm_interconnect_2_ocm_256k_dma_s2_chipselect;                      // mm_interconnect_2:ocm_256k_dma_s2_chipselect -> ocm_256k_dma:chipselect2
	wire   [63:0] mm_interconnect_2_ocm_256k_dma_s2_readdata;                        // ocm_256k_dma:readdata2 -> mm_interconnect_2:ocm_256k_dma_s2_readdata
	wire   [14:0] mm_interconnect_2_ocm_256k_dma_s2_address;                         // mm_interconnect_2:ocm_256k_dma_s2_address -> ocm_256k_dma:address2
	wire    [7:0] mm_interconnect_2_ocm_256k_dma_s2_byteenable;                      // mm_interconnect_2:ocm_256k_dma_s2_byteenable -> ocm_256k_dma:byteenable2
	wire          mm_interconnect_2_ocm_256k_dma_s2_write;                           // mm_interconnect_2:ocm_256k_dma_s2_write -> ocm_256k_dma:write2
	wire   [63:0] mm_interconnect_2_ocm_256k_dma_s2_writedata;                       // mm_interconnect_2:ocm_256k_dma_s2_writedata -> ocm_256k_dma:writedata2
	wire          mm_interconnect_2_ocm_256k_dma_s2_clken;                           // mm_interconnect_2:ocm_256k_dma_s2_clken -> ocm_256k_dma:clken2
	wire          mm_interconnect_2_pcie_256_dma_wr_dts_slave_chipselect;            // mm_interconnect_2:pcie_256_dma_wr_dts_slave_chipselect -> pcie_256_dma:WrDTSChipSelect_i
	wire          mm_interconnect_2_pcie_256_dma_wr_dts_slave_waitrequest;           // pcie_256_dma:WrDTSWaitRequest_o -> mm_interconnect_2:pcie_256_dma_wr_dts_slave_waitrequest
	wire    [7:0] mm_interconnect_2_pcie_256_dma_wr_dts_slave_address;               // mm_interconnect_2:pcie_256_dma_wr_dts_slave_address -> pcie_256_dma:WrDTSAddress_i
	wire          mm_interconnect_2_pcie_256_dma_wr_dts_slave_write;                 // mm_interconnect_2:pcie_256_dma_wr_dts_slave_write -> pcie_256_dma:WrDTSWrite_i
	wire  [255:0] mm_interconnect_2_pcie_256_dma_wr_dts_slave_writedata;             // mm_interconnect_2:pcie_256_dma_wr_dts_slave_writedata -> pcie_256_dma:WrDTSWriteData_i
	wire    [4:0] mm_interconnect_2_pcie_256_dma_wr_dts_slave_burstcount;            // mm_interconnect_2:pcie_256_dma_wr_dts_slave_burstcount -> pcie_256_dma:WrDTSBurstCount_i
	wire          alt_vip_cl_vfb_0_mem_master_rd_waitrequest;                        // mm_interconnect_3:alt_vip_cl_vfb_0_mem_master_rd_waitrequest -> alt_vip_cl_vfb_0:mem_master_rd_waitrequest
	wire   [31:0] alt_vip_cl_vfb_0_mem_master_rd_readdata;                           // mm_interconnect_3:alt_vip_cl_vfb_0_mem_master_rd_readdata -> alt_vip_cl_vfb_0:mem_master_rd_readdata
	wire   [31:0] alt_vip_cl_vfb_0_mem_master_rd_address;                            // alt_vip_cl_vfb_0:mem_master_rd_address -> mm_interconnect_3:alt_vip_cl_vfb_0_mem_master_rd_address
	wire          alt_vip_cl_vfb_0_mem_master_rd_read;                               // alt_vip_cl_vfb_0:mem_master_rd_read -> mm_interconnect_3:alt_vip_cl_vfb_0_mem_master_rd_read
	wire          alt_vip_cl_vfb_0_mem_master_rd_readdatavalid;                      // mm_interconnect_3:alt_vip_cl_vfb_0_mem_master_rd_readdatavalid -> alt_vip_cl_vfb_0:mem_master_rd_readdatavalid
	wire    [5:0] alt_vip_cl_vfb_0_mem_master_rd_burstcount;                         // alt_vip_cl_vfb_0:mem_master_rd_burstcount -> mm_interconnect_3:alt_vip_cl_vfb_0_mem_master_rd_burstcount
	wire          alt_vip_cl_vfb_0_mem_master_wr_waitrequest;                        // mm_interconnect_3:alt_vip_cl_vfb_0_mem_master_wr_waitrequest -> alt_vip_cl_vfb_0:mem_master_wr_waitrequest
	wire   [31:0] alt_vip_cl_vfb_0_mem_master_wr_address;                            // alt_vip_cl_vfb_0:mem_master_wr_address -> mm_interconnect_3:alt_vip_cl_vfb_0_mem_master_wr_address
	wire    [3:0] alt_vip_cl_vfb_0_mem_master_wr_byteenable;                         // alt_vip_cl_vfb_0:mem_master_wr_byteenable -> mm_interconnect_3:alt_vip_cl_vfb_0_mem_master_wr_byteenable
	wire          alt_vip_cl_vfb_0_mem_master_wr_write;                              // alt_vip_cl_vfb_0:mem_master_wr_write -> mm_interconnect_3:alt_vip_cl_vfb_0_mem_master_wr_write
	wire   [31:0] alt_vip_cl_vfb_0_mem_master_wr_writedata;                          // alt_vip_cl_vfb_0:mem_master_wr_writedata -> mm_interconnect_3:alt_vip_cl_vfb_0_mem_master_wr_writedata
	wire    [5:0] alt_vip_cl_vfb_0_mem_master_wr_burstcount;                         // alt_vip_cl_vfb_0:mem_master_wr_burstcount -> mm_interconnect_3:alt_vip_cl_vfb_0_mem_master_wr_burstcount
	wire          mm_interconnect_3_sdram_vfb_s1_chipselect;                         // mm_interconnect_3:sdram_vfb_s1_chipselect -> sdram_vfb:az_cs
	wire   [15:0] mm_interconnect_3_sdram_vfb_s1_readdata;                           // sdram_vfb:za_data -> mm_interconnect_3:sdram_vfb_s1_readdata
	wire          mm_interconnect_3_sdram_vfb_s1_waitrequest;                        // sdram_vfb:za_waitrequest -> mm_interconnect_3:sdram_vfb_s1_waitrequest
	wire   [24:0] mm_interconnect_3_sdram_vfb_s1_address;                            // mm_interconnect_3:sdram_vfb_s1_address -> sdram_vfb:az_addr
	wire          mm_interconnect_3_sdram_vfb_s1_read;                               // mm_interconnect_3:sdram_vfb_s1_read -> sdram_vfb:az_rd_n
	wire    [1:0] mm_interconnect_3_sdram_vfb_s1_byteenable;                         // mm_interconnect_3:sdram_vfb_s1_byteenable -> sdram_vfb:az_be_n
	wire          mm_interconnect_3_sdram_vfb_s1_readdatavalid;                      // sdram_vfb:za_valid -> mm_interconnect_3:sdram_vfb_s1_readdatavalid
	wire          mm_interconnect_3_sdram_vfb_s1_write;                              // mm_interconnect_3:sdram_vfb_s1_write -> sdram_vfb:az_wr_n
	wire   [15:0] mm_interconnect_3_sdram_vfb_s1_writedata;                          // mm_interconnect_3:sdram_vfb_s1_writedata -> sdram_vfb:az_data
	wire          pcie_256_dma_rd_dcm_master_waitrequest;                            // mm_interconnect_4:pcie_256_dma_rd_dcm_master_waitrequest -> pcie_256_dma:RdDCMWaitRequest_i
	wire   [31:0] pcie_256_dma_rd_dcm_master_readdata;                               // mm_interconnect_4:pcie_256_dma_rd_dcm_master_readdata -> pcie_256_dma:RdDCMReadData_i
	wire   [63:0] pcie_256_dma_rd_dcm_master_address;                                // pcie_256_dma:RdDCMAddress_o -> mm_interconnect_4:pcie_256_dma_rd_dcm_master_address
	wire          pcie_256_dma_rd_dcm_master_read;                                   // pcie_256_dma:RdDCMRead_o -> mm_interconnect_4:pcie_256_dma_rd_dcm_master_read
	wire    [3:0] pcie_256_dma_rd_dcm_master_byteenable;                             // pcie_256_dma:RdDCMByteEnable_o -> mm_interconnect_4:pcie_256_dma_rd_dcm_master_byteenable
	wire          pcie_256_dma_rd_dcm_master_readdatavalid;                          // mm_interconnect_4:pcie_256_dma_rd_dcm_master_readdatavalid -> pcie_256_dma:RdDCMReadDataValid_i
	wire          pcie_256_dma_rd_dcm_master_write;                                  // pcie_256_dma:RdDCMWrite_o -> mm_interconnect_4:pcie_256_dma_rd_dcm_master_write
	wire   [31:0] pcie_256_dma_rd_dcm_master_writedata;                              // pcie_256_dma:RdDCMWriteData_o -> mm_interconnect_4:pcie_256_dma_rd_dcm_master_writedata
	wire          pcie_256_dma_wr_dcm_master_waitrequest;                            // mm_interconnect_4:pcie_256_dma_wr_dcm_master_waitrequest -> pcie_256_dma:WrDCMWaitRequest_i
	wire   [31:0] pcie_256_dma_wr_dcm_master_readdata;                               // mm_interconnect_4:pcie_256_dma_wr_dcm_master_readdata -> pcie_256_dma:WrDCMReadData_i
	wire   [63:0] pcie_256_dma_wr_dcm_master_address;                                // pcie_256_dma:WrDCMAddress_o -> mm_interconnect_4:pcie_256_dma_wr_dcm_master_address
	wire          pcie_256_dma_wr_dcm_master_read;                                   // pcie_256_dma:WrDCMRead_o -> mm_interconnect_4:pcie_256_dma_wr_dcm_master_read
	wire    [3:0] pcie_256_dma_wr_dcm_master_byteenable;                             // pcie_256_dma:WrDCMByteEnable_o -> mm_interconnect_4:pcie_256_dma_wr_dcm_master_byteenable
	wire          pcie_256_dma_wr_dcm_master_readdatavalid;                          // mm_interconnect_4:pcie_256_dma_wr_dcm_master_readdatavalid -> pcie_256_dma:WrDCMReadDataValid_i
	wire          pcie_256_dma_wr_dcm_master_write;                                  // pcie_256_dma:WrDCMWrite_o -> mm_interconnect_4:pcie_256_dma_wr_dcm_master_write
	wire   [31:0] pcie_256_dma_wr_dcm_master_writedata;                              // pcie_256_dma:WrDCMWriteData_o -> mm_interconnect_4:pcie_256_dma_wr_dcm_master_writedata
	wire          mm_interconnect_4_pcie_256_dma_txs_chipselect;                     // mm_interconnect_4:pcie_256_dma_Txs_chipselect -> pcie_256_dma:TxsChipSelect_i
	wire   [31:0] mm_interconnect_4_pcie_256_dma_txs_readdata;                       // pcie_256_dma:TxsReadData_o -> mm_interconnect_4:pcie_256_dma_Txs_readdata
	wire          mm_interconnect_4_pcie_256_dma_txs_waitrequest;                    // pcie_256_dma:TxsWaitRequest_o -> mm_interconnect_4:pcie_256_dma_Txs_waitrequest
	wire   [63:0] mm_interconnect_4_pcie_256_dma_txs_address;                        // mm_interconnect_4:pcie_256_dma_Txs_address -> pcie_256_dma:TxsAddress_i
	wire          mm_interconnect_4_pcie_256_dma_txs_read;                           // mm_interconnect_4:pcie_256_dma_Txs_read -> pcie_256_dma:TxsRead_i
	wire    [3:0] mm_interconnect_4_pcie_256_dma_txs_byteenable;                     // mm_interconnect_4:pcie_256_dma_Txs_byteenable -> pcie_256_dma:TxsByteEnable_i
	wire          mm_interconnect_4_pcie_256_dma_txs_readdatavalid;                  // pcie_256_dma:TxsReadDataValid_o -> mm_interconnect_4:pcie_256_dma_Txs_readdatavalid
	wire          mm_interconnect_4_pcie_256_dma_txs_write;                          // mm_interconnect_4:pcie_256_dma_Txs_write -> pcie_256_dma:TxsWrite_i
	wire   [31:0] mm_interconnect_4_pcie_256_dma_txs_writedata;                      // mm_interconnect_4:pcie_256_dma_Txs_writedata -> pcie_256_dma:TxsWriteData_i
	wire   [31:0] pcie_reconfig_driver_0_reconfig_mgmt_readdata;                     // mm_interconnect_5:pcie_reconfig_driver_0_reconfig_mgmt_readdata -> pcie_reconfig_driver_0:reconfig_mgmt_readdata
	wire          pcie_reconfig_driver_0_reconfig_mgmt_waitrequest;                  // mm_interconnect_5:pcie_reconfig_driver_0_reconfig_mgmt_waitrequest -> pcie_reconfig_driver_0:reconfig_mgmt_waitrequest
	wire    [6:0] pcie_reconfig_driver_0_reconfig_mgmt_address;                      // pcie_reconfig_driver_0:reconfig_mgmt_address -> mm_interconnect_5:pcie_reconfig_driver_0_reconfig_mgmt_address
	wire          pcie_reconfig_driver_0_reconfig_mgmt_read;                         // pcie_reconfig_driver_0:reconfig_mgmt_read -> mm_interconnect_5:pcie_reconfig_driver_0_reconfig_mgmt_read
	wire          pcie_reconfig_driver_0_reconfig_mgmt_write;                        // pcie_reconfig_driver_0:reconfig_mgmt_write -> mm_interconnect_5:pcie_reconfig_driver_0_reconfig_mgmt_write
	wire   [31:0] pcie_reconfig_driver_0_reconfig_mgmt_writedata;                    // pcie_reconfig_driver_0:reconfig_mgmt_writedata -> mm_interconnect_5:pcie_reconfig_driver_0_reconfig_mgmt_writedata
	wire   [31:0] mm_interconnect_5_alt_xcvr_reconfig_0_reconfig_mgmt_readdata;      // alt_xcvr_reconfig_0:reconfig_mgmt_readdata -> mm_interconnect_5:alt_xcvr_reconfig_0_reconfig_mgmt_readdata
	wire          mm_interconnect_5_alt_xcvr_reconfig_0_reconfig_mgmt_waitrequest;   // alt_xcvr_reconfig_0:reconfig_mgmt_waitrequest -> mm_interconnect_5:alt_xcvr_reconfig_0_reconfig_mgmt_waitrequest
	wire    [6:0] mm_interconnect_5_alt_xcvr_reconfig_0_reconfig_mgmt_address;       // mm_interconnect_5:alt_xcvr_reconfig_0_reconfig_mgmt_address -> alt_xcvr_reconfig_0:reconfig_mgmt_address
	wire          mm_interconnect_5_alt_xcvr_reconfig_0_reconfig_mgmt_read;          // mm_interconnect_5:alt_xcvr_reconfig_0_reconfig_mgmt_read -> alt_xcvr_reconfig_0:reconfig_mgmt_read
	wire          mm_interconnect_5_alt_xcvr_reconfig_0_reconfig_mgmt_write;         // mm_interconnect_5:alt_xcvr_reconfig_0_reconfig_mgmt_write -> alt_xcvr_reconfig_0:reconfig_mgmt_write
	wire   [31:0] mm_interconnect_5_alt_xcvr_reconfig_0_reconfig_mgmt_writedata;     // mm_interconnect_5:alt_xcvr_reconfig_0_reconfig_mgmt_writedata -> alt_xcvr_reconfig_0:reconfig_mgmt_writedata
	wire          irq_mapper_receiver0_irq;                                          // fifo_0:wrclk_control_slave_irq -> irq_mapper:receiver0_irq
	wire          irq_mapper_receiver1_irq;                                          // i2c_opencores_mipi:wb_inta_o -> irq_mapper:receiver1_irq
	wire          irq_mapper_receiver2_irq;                                          // i2c_opencores_camera:wb_inta_o -> irq_mapper:receiver2_irq
	wire          irq_mapper_receiver3_irq;                                          // jtag_uart_0:av_irq -> irq_mapper:receiver3_irq
	wire          irq_mapper_receiver4_irq;                                          // pio_button:irq -> irq_mapper:receiver4_irq
	wire          irq_mapper_receiver5_irq;                                          // timer_0:irq -> irq_mapper:receiver5_irq
	wire   [31:0] nios2_gen2_0_irq_irq;                                              // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire          terasic_camera_0_avalon_streaming_source_valid;                    // TERASIC_CAMERA_0:st_valid -> avalon_st_adapter:in_0_valid
	wire   [23:0] terasic_camera_0_avalon_streaming_source_data;                     // TERASIC_CAMERA_0:st_data -> avalon_st_adapter:in_0_data
	wire          terasic_camera_0_avalon_streaming_source_ready;                    // avalon_st_adapter:in_0_ready -> TERASIC_CAMERA_0:st_ready
	wire          terasic_camera_0_avalon_streaming_source_startofpacket;            // TERASIC_CAMERA_0:st_sop -> avalon_st_adapter:in_0_startofpacket
	wire          terasic_camera_0_avalon_streaming_source_endofpacket;              // TERASIC_CAMERA_0:st_eop -> avalon_st_adapter:in_0_endofpacket
	wire          avalon_st_adapter_out_0_valid;                                     // avalon_st_adapter:out_0_valid -> alt_vip_cl_vfb_0:din_valid
	wire   [23:0] avalon_st_adapter_out_0_data;                                      // avalon_st_adapter:out_0_data -> alt_vip_cl_vfb_0:din_data
	wire          avalon_st_adapter_out_0_ready;                                     // alt_vip_cl_vfb_0:din_ready -> avalon_st_adapter:out_0_ready
	wire          avalon_st_adapter_out_0_startofpacket;                             // avalon_st_adapter:out_0_startofpacket -> alt_vip_cl_vfb_0:din_startofpacket
	wire          avalon_st_adapter_out_0_endofpacket;                               // avalon_st_adapter:out_0_endofpacket -> alt_vip_cl_vfb_0:din_endofpacket
	wire          terasic_auto_focus_0_dout_valid;                                   // TERASIC_AUTO_FOCUS_0:source_valid -> avalon_st_adapter_001:in_0_valid
	wire   [31:0] terasic_auto_focus_0_dout_data;                                    // TERASIC_AUTO_FOCUS_0:source_data -> avalon_st_adapter_001:in_0_data
	wire          terasic_auto_focus_0_dout_ready;                                   // avalon_st_adapter_001:in_0_ready -> TERASIC_AUTO_FOCUS_0:source_ready
	wire          terasic_auto_focus_0_dout_startofpacket;                           // TERASIC_AUTO_FOCUS_0:source_sop -> avalon_st_adapter_001:in_0_startofpacket
	wire          terasic_auto_focus_0_dout_endofpacket;                             // TERASIC_AUTO_FOCUS_0:source_eop -> avalon_st_adapter_001:in_0_endofpacket
	wire          avalon_st_adapter_001_out_0_valid;                                 // avalon_st_adapter_001:out_0_valid -> fifo_0:avalonst_sink_valid
	wire   [31:0] avalon_st_adapter_001_out_0_data;                                  // avalon_st_adapter_001:out_0_data -> fifo_0:avalonst_sink_data
	wire          avalon_st_adapter_001_out_0_ready;                                 // fifo_0:avalonst_sink_ready -> avalon_st_adapter_001:out_0_ready
	wire    [7:0] avalon_st_adapter_001_out_0_channel;                               // avalon_st_adapter_001:out_0_channel -> fifo_0:avalonst_sink_channel
	wire          avalon_st_adapter_001_out_0_startofpacket;                         // avalon_st_adapter_001:out_0_startofpacket -> fifo_0:avalonst_sink_startofpacket
	wire          avalon_st_adapter_001_out_0_endofpacket;                           // avalon_st_adapter_001:out_0_endofpacket -> fifo_0:avalonst_sink_endofpacket
	wire    [7:0] avalon_st_adapter_001_out_0_error;                                 // avalon_st_adapter_001:out_0_error -> fifo_0:avalonst_sink_error
	wire    [1:0] avalon_st_adapter_001_out_0_empty;                                 // avalon_st_adapter_001:out_0_empty -> fifo_0:avalonst_sink_empty
	wire          rst_controller_reset_out_reset;                                    // rst_controller:reset_out -> [TERASIC_AUTO_FOCUS_0:reset_n, TERASIC_CAMERA_0:reset_n, alt_vip_cl_vfb_0:main_reset, avalon_st_adapter:in_rst_0_reset, avalon_st_adapter_001:in_rst_0_reset, csr_regmap:reset, ddr3_status:reset_n, fifo_0:reset_n, i2c_opencores_camera:wb_rst_i, i2c_opencores_mipi:wb_rst_i, irq_mapper:reset, jtag_uart_0:rst_n, mipi_pwdn_n:reset_n, mipi_reset_n:reset_n, mm_interconnect_1:mem_if_ddr3_emif_0_mp_cmd_reset_n_0_reset_bridge_in_reset_reset, mm_interconnect_1:nios2_gen2_0_reset_reset_bridge_in_reset_reset, mm_interconnect_3:alt_vip_cl_vfb_0_main_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, nios_ram:reset, ocm_256k_dma:reset, pio_button:reset_n, pio_led:reset_n, rst_translator:in_reset, sdram_vfb:reset_n, sysid_qsys_0:reset_n, timer_0:reset_n]
	wire          rst_controller_reset_out_reset_req;                                // rst_controller:reset_req -> [csr_regmap:reset_req, nios2_gen2_0:reset_req, nios_ram:reset_req, ocm_256k_dma:reset_req, rst_translator:reset_req_in]
	wire          rst_controller_001_reset_out_reset;                                // rst_controller_001:reset_out -> [alt_xcvr_reconfig_0:mgmt_rst_reset, mm_interconnect_5:alt_xcvr_reconfig_0_mgmt_rst_reset_reset_bridge_in_reset_reset]
	wire          rst_controller_002_reset_out_reset;                                // rst_controller_002:reset_out -> [csr_regmap:reset2, mm_interconnect_0:csr_regmap_reset2_reset_bridge_in_reset_reset, mm_interconnect_2:ocm_256k_dma_reset2_reset_bridge_in_reset_reset, mm_interconnect_4:pcie_256_dma_rd_dcm_master_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_5:pcie_reconfig_driver_0_reconfig_xcvr_rst_reset_bridge_in_reset_reset, ocm_256k_dma:reset2, pcie_reconfig_driver_0:reconfig_xcvr_rst, rst_translator_001:in_reset]
	wire          rst_controller_002_reset_out_reset_req;                            // rst_controller_002:reset_req -> [csr_regmap:reset_req2, ocm_256k_dma:reset_req2, rst_translator_001:reset_req_in]
	wire          pcie_256_dma_nreset_status_reset;                                  // pcie_256_dma:reset_status -> rst_controller_002:reset_in0

	TERASIC_AUTO_FOCUS #(
		.VIDEO_W (640),
		.VIDEO_H (480)
	) terasic_auto_focus_0 (
		.clk          (pll_0_outclk0_clk),                                         //   clock.clk
		.reset_n      (~rst_controller_reset_out_reset),                           //   reset.reset_n
		.s_chipselect (mm_interconnect_1_terasic_auto_focus_0_mm_ctrl_chipselect), // mm_ctrl.chipselect
		.s_read       (mm_interconnect_1_terasic_auto_focus_0_mm_ctrl_read),       //        .read
		.s_write      (mm_interconnect_1_terasic_auto_focus_0_mm_ctrl_write),      //        .write
		.s_readdata   (mm_interconnect_1_terasic_auto_focus_0_mm_ctrl_readdata),   //        .readdata
		.s_writedata  (mm_interconnect_1_terasic_auto_focus_0_mm_ctrl_writedata),  //        .writedata
		.s_address    (mm_interconnect_1_terasic_auto_focus_0_mm_ctrl_address),    //        .address
		.sink_data    (alt_vip_cl_vfb_0_dout_data),                                //     din.data
		.sink_valid   (alt_vip_cl_vfb_0_dout_valid),                               //        .valid
		.sink_ready   (alt_vip_cl_vfb_0_dout_ready),                               //        .ready
		.sink_sop     (alt_vip_cl_vfb_0_dout_startofpacket),                       //        .startofpacket
		.sink_eop     (alt_vip_cl_vfb_0_dout_endofpacket),                         //        .endofpacket
		.source_data  (terasic_auto_focus_0_dout_data),                            //    dout.data
		.source_valid (terasic_auto_focus_0_dout_valid),                           //        .valid
		.source_ready (terasic_auto_focus_0_dout_ready),                           //        .ready
		.source_sop   (terasic_auto_focus_0_dout_startofpacket),                   //        .startofpacket
		.source_eop   (terasic_auto_focus_0_dout_endofpacket),                     //        .endofpacket
		.vcm_i2c_sda  (terasic_auto_focus_0_conduit_vcm_i2c_sda),                  // Conduit.vcm_i2c_sda
		.clk50        (terasic_auto_focus_0_conduit_clk50),                        //        .clk50
		.vcm_i2c_scl  (terasic_auto_focus_0_conduit_vcm_i2c_scl)                   //        .vcm_i2c_scl
	);

	TERASIC_CAMERA #(
		.VIDEO_W (640),
		.VIDEO_H (480)
	) terasic_camera_0 (
		.clk           (pll_0_outclk0_clk),                                      //             clock_reset.clk
		.reset_n       (~rst_controller_reset_out_reset),                        //       clock_reset_reset.reset_n
		.CAMERA_D      (terasic_camera_0_conduit_end_cam_d),                     //             conduit_end.cam_d
		.CAMERA_FVAL   (terasic_camera_0_conduit_end_cam_fval),                  //                        .cam_fval
		.CAMERA_LVAL   (terasic_camera_0_conduit_end_cam_lval),                  //                        .cam_lval
		.CAMERA_PIXCLK (terasic_camera_0_conduit_end_cam_pix),                   //                        .cam_pix
		.st_data       (terasic_camera_0_avalon_streaming_source_data),          // avalon_streaming_source.data
		.st_valid      (terasic_camera_0_avalon_streaming_source_valid),         //                        .valid
		.st_sop        (terasic_camera_0_avalon_streaming_source_startofpacket), //                        .startofpacket
		.st_eop        (terasic_camera_0_avalon_streaming_source_endofpacket),   //                        .endofpacket
		.st_ready      (terasic_camera_0_avalon_streaming_source_ready)          //                        .ready
	);

	top_alt_vip_cl_vfb_0 #(
		.BITS_PER_SYMBOL              (8),
		.NUMBER_OF_COLOR_PLANES       (3),
		.COLOR_PLANES_ARE_IN_PARALLEL (1),
		.PIXELS_IN_PARALLEL           (1),
		.READY_LATENCY                (1),
		.MAX_WIDTH                    (640),
		.MAX_HEIGHT                   (480),
		.CLOCKS_ARE_SEPARATE          (0),
		.MEM_PORT_WIDTH               (32),
		.MEM_BASE_ADDR                (0),
		.BURST_ALIGNMENT              (1),
		.WRITE_FIFO_DEPTH             (512),
		.WRITE_BURST_TARGET           (32),
		.READ_FIFO_DEPTH              (512),
		.READ_BURST_TARGET            (32),
		.WRITER_RUNTIME_CONTROL       (0),
		.READER_RUNTIME_CONTROL       (0),
		.IS_FRAME_WRITER              (0),
		.IS_FRAME_READER              (0),
		.DROP_FRAMES                  (1),
		.REPEAT_FRAMES                (1),
		.DROP_REPEAT_USER             (0),
		.INTERLACED_SUPPORT           (0),
		.CONTROLLED_DROP_REPEAT       (0),
		.DROP_INVALID_FIELDS          (0),
		.MULTI_FRAME_DELAY            (1),
		.IS_SYNC_MASTER               (0),
		.IS_SYNC_SLAVE                (0),
		.LINE_BASED_BUFFERING         (0),
		.PRIORITIZE_FMAX              (0),
		.USER_PACKETS_MAX_STORAGE     (1),
		.MAX_SYMBOLS_PER_PACKET       (10),
		.NUM_BUFFERS                  (3)
	) alt_vip_cl_vfb_0 (
		.main_clock                  (pll_0_outclk0_clk),                            //    main_clock.clk
		.main_reset                  (rst_controller_reset_out_reset),               //    main_reset.reset
		.din_data                    (avalon_st_adapter_out_0_data),                 //           din.data
		.din_valid                   (avalon_st_adapter_out_0_valid),                //              .valid
		.din_startofpacket           (avalon_st_adapter_out_0_startofpacket),        //              .startofpacket
		.din_endofpacket             (avalon_st_adapter_out_0_endofpacket),          //              .endofpacket
		.din_ready                   (avalon_st_adapter_out_0_ready),                //              .ready
		.mem_master_wr_address       (alt_vip_cl_vfb_0_mem_master_wr_address),       // mem_master_wr.address
		.mem_master_wr_burstcount    (alt_vip_cl_vfb_0_mem_master_wr_burstcount),    //              .burstcount
		.mem_master_wr_waitrequest   (alt_vip_cl_vfb_0_mem_master_wr_waitrequest),   //              .waitrequest
		.mem_master_wr_write         (alt_vip_cl_vfb_0_mem_master_wr_write),         //              .write
		.mem_master_wr_writedata     (alt_vip_cl_vfb_0_mem_master_wr_writedata),     //              .writedata
		.mem_master_wr_byteenable    (alt_vip_cl_vfb_0_mem_master_wr_byteenable),    //              .byteenable
		.dout_data                   (alt_vip_cl_vfb_0_dout_data),                   //          dout.data
		.dout_valid                  (alt_vip_cl_vfb_0_dout_valid),                  //              .valid
		.dout_startofpacket          (alt_vip_cl_vfb_0_dout_startofpacket),          //              .startofpacket
		.dout_endofpacket            (alt_vip_cl_vfb_0_dout_endofpacket),            //              .endofpacket
		.dout_ready                  (alt_vip_cl_vfb_0_dout_ready),                  //              .ready
		.mem_master_rd_address       (alt_vip_cl_vfb_0_mem_master_rd_address),       // mem_master_rd.address
		.mem_master_rd_burstcount    (alt_vip_cl_vfb_0_mem_master_rd_burstcount),    //              .burstcount
		.mem_master_rd_waitrequest   (alt_vip_cl_vfb_0_mem_master_rd_waitrequest),   //              .waitrequest
		.mem_master_rd_read          (alt_vip_cl_vfb_0_mem_master_rd_read),          //              .read
		.mem_master_rd_readdata      (alt_vip_cl_vfb_0_mem_master_rd_readdata),      //              .readdata
		.mem_master_rd_readdatavalid (alt_vip_cl_vfb_0_mem_master_rd_readdatavalid)  //              .readdatavalid
	);

	alt_xcvr_reconfig #(
		.device_family                 ("Cyclone V"),
		.number_of_reconfig_interfaces (5),
		.enable_offset                 (1),
		.enable_lc                     (0),
		.enable_dcd                    (0),
		.enable_dcd_power_up           (1),
		.enable_analog                 (1),
		.enable_eyemon                 (0),
		.enable_ber                    (0),
		.enable_dfe                    (0),
		.enable_adce                   (1),
		.enable_mif                    (0),
		.enable_pll                    (0)
	) alt_xcvr_reconfig_0 (
		.reconfig_busy             (),                                                                //      reconfig_busy.reconfig_busy
		.mgmt_clk_clk              (clk_clk),                                                         //       mgmt_clk_clk.clk
		.mgmt_rst_reset            (rst_controller_001_reset_out_reset),                              //     mgmt_rst_reset.reset
		.reconfig_mgmt_address     (mm_interconnect_5_alt_xcvr_reconfig_0_reconfig_mgmt_address),     //      reconfig_mgmt.address
		.reconfig_mgmt_read        (mm_interconnect_5_alt_xcvr_reconfig_0_reconfig_mgmt_read),        //                   .read
		.reconfig_mgmt_readdata    (mm_interconnect_5_alt_xcvr_reconfig_0_reconfig_mgmt_readdata),    //                   .readdata
		.reconfig_mgmt_waitrequest (mm_interconnect_5_alt_xcvr_reconfig_0_reconfig_mgmt_waitrequest), //                   .waitrequest
		.reconfig_mgmt_write       (mm_interconnect_5_alt_xcvr_reconfig_0_reconfig_mgmt_write),       //                   .write
		.reconfig_mgmt_writedata   (mm_interconnect_5_alt_xcvr_reconfig_0_reconfig_mgmt_writedata),   //                   .writedata
		.reconfig_to_xcvr          (alt_xcvr_reconfig_0_reconfig_to_xcvr_reconfig_to_xcvr),           //   reconfig_to_xcvr.reconfig_to_xcvr
		.reconfig_from_xcvr        (pcie_256_dma_reconfig_from_xcvr_reconfig_from_xcvr),              // reconfig_from_xcvr.reconfig_from_xcvr
		.tx_cal_busy               (),                                                                //        (terminated)
		.rx_cal_busy               (),                                                                //        (terminated)
		.cal_busy_in               (1'b0),                                                            //        (terminated)
		.reconfig_mif_address      (),                                                                //        (terminated)
		.reconfig_mif_read         (),                                                                //        (terminated)
		.reconfig_mif_readdata     (16'b0000000000000000),                                            //        (terminated)
		.reconfig_mif_waitrequest  (1'b0)                                                             //        (terminated)
	);

	top_csr_regmap csr_regmap (
		.clk         (pll_0_outclk0_clk),                          //   clk1.clk
		.address     (mm_interconnect_1_csr_regmap_s1_address),    //     s1.address
		.clken       (mm_interconnect_1_csr_regmap_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_1_csr_regmap_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_1_csr_regmap_s1_write),      //       .write
		.readdata    (mm_interconnect_1_csr_regmap_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_1_csr_regmap_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_1_csr_regmap_s1_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),             // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),         //       .reset_req
		.address2    (mm_interconnect_0_csr_regmap_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_0_csr_regmap_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_0_csr_regmap_s2_clken),      //       .clken
		.write2      (mm_interconnect_0_csr_regmap_s2_write),      //       .write
		.readdata2   (mm_interconnect_0_csr_regmap_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_0_csr_regmap_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_0_csr_regmap_s2_byteenable), //       .byteenable
		.clk2        (pcie_256_dma_coreclkout_clk),                //   clk2.clk
		.reset2      (rst_controller_002_reset_out_reset),         // reset2.reset
		.reset_req2  (rst_controller_002_reset_out_reset_req),     //       .reset_req
		.freeze      (1'b0)                                        // (terminated)
	);

	top_ddr3_status ddr3_status (
		.clk      (pll_0_outclk0_clk),                         //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_1_ddr3_status_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_ddr3_status_s1_readdata), //                    .readdata
		.in_port  (ddr3_status_external_connection_export)     // external_connection.export
	);

	top_fifo_0 fifo_0 (
		.wrclock                         (pll_0_outclk0_clk),                         //   clk_in.clk
		.reset_n                         (~rst_controller_reset_out_reset),           // reset_in.reset_n
		.avalonst_sink_valid             (avalon_st_adapter_001_out_0_valid),         //       in.valid
		.avalonst_sink_data              (avalon_st_adapter_001_out_0_data),          //         .data
		.avalonst_sink_channel           (avalon_st_adapter_001_out_0_channel),       //         .channel
		.avalonst_sink_error             (avalon_st_adapter_001_out_0_error),         //         .error
		.avalonst_sink_startofpacket     (avalon_st_adapter_001_out_0_startofpacket), //         .startofpacket
		.avalonst_sink_endofpacket       (avalon_st_adapter_001_out_0_endofpacket),   //         .endofpacket
		.avalonst_sink_empty             (avalon_st_adapter_001_out_0_empty),         //         .empty
		.avalonst_sink_ready             (avalon_st_adapter_001_out_0_ready),         //         .ready
		.avalonmm_read_slave_readdata    (mm_interconnect_1_fifo_0_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read        (mm_interconnect_1_fifo_0_out_read),         //         .read
		.avalonmm_read_slave_address     (mm_interconnect_1_fifo_0_out_address),      //         .address
		.avalonmm_read_slave_waitrequest (mm_interconnect_1_fifo_0_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address     (mm_interconnect_1_fifo_0_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read        (mm_interconnect_1_fifo_0_in_csr_read),      //         .read
		.wrclk_control_slave_writedata   (mm_interconnect_1_fifo_0_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write       (mm_interconnect_1_fifo_0_in_csr_write),     //         .write
		.wrclk_control_slave_readdata    (mm_interconnect_1_fifo_0_in_csr_readdata),  //         .readdata
		.wrclk_control_slave_irq         (irq_mapper_receiver0_irq)                   //   in_irq.irq
	);

	i2c_opencores i2c_opencores_camera (
		.wb_clk_i   (pll_0_outclk0_clk),                                                 //            clock.clk
		.wb_rst_i   (rst_controller_reset_out_reset),                                    //      clock_reset.reset
		.scl_pad_io (i2c_opencores_camera_export_scl_pad_io),                            //           export.scl_pad_io
		.sda_pad_io (i2c_opencores_camera_export_sda_pad_io),                            //                 .sda_pad_io
		.wb_adr_i   (mm_interconnect_1_i2c_opencores_camera_avalon_slave_0_address),     //   avalon_slave_0.address
		.wb_dat_i   (mm_interconnect_1_i2c_opencores_camera_avalon_slave_0_writedata),   //                 .writedata
		.wb_dat_o   (mm_interconnect_1_i2c_opencores_camera_avalon_slave_0_readdata),    //                 .readdata
		.wb_we_i    (mm_interconnect_1_i2c_opencores_camera_avalon_slave_0_write),       //                 .write
		.wb_stb_i   (mm_interconnect_1_i2c_opencores_camera_avalon_slave_0_chipselect),  //                 .chipselect
		.wb_ack_o   (mm_interconnect_1_i2c_opencores_camera_avalon_slave_0_waitrequest), //                 .waitrequest_n
		.wb_inta_o  (irq_mapper_receiver2_irq)                                           // interrupt_sender.irq
	);

	i2c_opencores i2c_opencores_mipi (
		.wb_clk_i   (pll_0_outclk0_clk),                                               //            clock.clk
		.wb_rst_i   (rst_controller_reset_out_reset),                                  //      clock_reset.reset
		.scl_pad_io (i2c_opencores_mipi_export_scl_pad_io),                            //           export.scl_pad_io
		.sda_pad_io (i2c_opencores_mipi_export_sda_pad_io),                            //                 .sda_pad_io
		.wb_adr_i   (mm_interconnect_1_i2c_opencores_mipi_avalon_slave_0_address),     //   avalon_slave_0.address
		.wb_dat_i   (mm_interconnect_1_i2c_opencores_mipi_avalon_slave_0_writedata),   //                 .writedata
		.wb_dat_o   (mm_interconnect_1_i2c_opencores_mipi_avalon_slave_0_readdata),    //                 .readdata
		.wb_we_i    (mm_interconnect_1_i2c_opencores_mipi_avalon_slave_0_write),       //                 .write
		.wb_stb_i   (mm_interconnect_1_i2c_opencores_mipi_avalon_slave_0_chipselect),  //                 .chipselect
		.wb_ack_o   (mm_interconnect_1_i2c_opencores_mipi_avalon_slave_0_waitrequest), //                 .waitrequest_n
		.wb_inta_o  (irq_mapper_receiver1_irq)                                         // interrupt_sender.irq
	);

	top_jtag_uart_0 jtag_uart_0 (
		.clk            (pll_0_outclk0_clk),                                           //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver3_irq)                                     //               irq.irq
	);

	top_mem_if_ddr3_emif_0 mem_if_ddr3_emif_0 (
		.pll_ref_clk                (mem_if_ddr3_emif_0_pll_ref_clk_clk),                            //        pll_ref_clk.clk
		.global_reset_n             (reset_reset_n),                                                 //       global_reset.reset_n
		.soft_reset_n               (reset_reset_n),                                                 //         soft_reset.reset_n
		.afi_clk                    (),                                                              //            afi_clk.clk
		.afi_half_clk               (),                                                              //       afi_half_clk.clk
		.afi_reset_n                (),                                                              //          afi_reset.reset_n
		.afi_reset_export_n         (),                                                              //   afi_reset_export.reset_n
		.mem_a                      (memory_mem_a),                                                  //             memory.mem_a
		.mem_ba                     (memory_mem_ba),                                                 //                   .mem_ba
		.mem_ck                     (memory_mem_ck),                                                 //                   .mem_ck
		.mem_ck_n                   (memory_mem_ck_n),                                               //                   .mem_ck_n
		.mem_cke                    (memory_mem_cke),                                                //                   .mem_cke
		.mem_cs_n                   (memory_mem_cs_n),                                               //                   .mem_cs_n
		.mem_dm                     (memory_mem_dm),                                                 //                   .mem_dm
		.mem_ras_n                  (memory_mem_ras_n),                                              //                   .mem_ras_n
		.mem_cas_n                  (memory_mem_cas_n),                                              //                   .mem_cas_n
		.mem_we_n                   (memory_mem_we_n),                                               //                   .mem_we_n
		.mem_reset_n                (memory_mem_reset_n),                                            //                   .mem_reset_n
		.mem_dq                     (memory_mem_dq),                                                 //                   .mem_dq
		.mem_dqs                    (memory_mem_dqs),                                                //                   .mem_dqs
		.mem_dqs_n                  (memory_mem_dqs_n),                                              //                   .mem_dqs_n
		.mem_odt                    (memory_mem_odt),                                                //                   .mem_odt
		.avl_ready_0                (mm_interconnect_1_mem_if_ddr3_emif_0_avl_0_waitrequest),        //              avl_0.waitrequest_n
		.avl_burstbegin_0           (mm_interconnect_1_mem_if_ddr3_emif_0_avl_0_beginbursttransfer), //                   .beginbursttransfer
		.avl_addr_0                 (mm_interconnect_1_mem_if_ddr3_emif_0_avl_0_address),            //                   .address
		.avl_rdata_valid_0          (mm_interconnect_1_mem_if_ddr3_emif_0_avl_0_readdatavalid),      //                   .readdatavalid
		.avl_rdata_0                (mm_interconnect_1_mem_if_ddr3_emif_0_avl_0_readdata),           //                   .readdata
		.avl_wdata_0                (mm_interconnect_1_mem_if_ddr3_emif_0_avl_0_writedata),          //                   .writedata
		.avl_be_0                   (mm_interconnect_1_mem_if_ddr3_emif_0_avl_0_byteenable),         //                   .byteenable
		.avl_read_req_0             (mm_interconnect_1_mem_if_ddr3_emif_0_avl_0_read),               //                   .read
		.avl_write_req_0            (mm_interconnect_1_mem_if_ddr3_emif_0_avl_0_write),              //                   .write
		.avl_size_0                 (mm_interconnect_1_mem_if_ddr3_emif_0_avl_0_burstcount),         //                   .burstcount
		.mp_cmd_clk_0_clk           (pll_0_outclk0_clk),                                             //       mp_cmd_clk_0.clk
		.mp_cmd_reset_n_0_reset_n   (reset_reset_n),                                                 //   mp_cmd_reset_n_0.reset_n
		.mp_rfifo_clk_0_clk         (pll_0_outclk0_clk),                                             //     mp_rfifo_clk_0.clk
		.mp_rfifo_reset_n_0_reset_n (reset_reset_n),                                                 // mp_rfifo_reset_n_0.reset_n
		.mp_wfifo_clk_0_clk         (pll_0_outclk0_clk),                                             //     mp_wfifo_clk_0.clk
		.mp_wfifo_reset_n_0_reset_n (reset_reset_n),                                                 // mp_wfifo_reset_n_0.reset_n
		.mp_rfifo_clk_1_clk         (pll_0_outclk0_clk),                                             //     mp_rfifo_clk_1.clk
		.mp_rfifo_reset_n_1_reset_n (reset_reset_n),                                                 // mp_rfifo_reset_n_1.reset_n
		.mp_wfifo_clk_1_clk         (pll_0_outclk0_clk),                                             //     mp_wfifo_clk_1.clk
		.mp_wfifo_reset_n_1_reset_n (reset_reset_n),                                                 // mp_wfifo_reset_n_1.reset_n
		.local_init_done            (mem_if_ddr3_emif_0_status_local_init_done),                     //             status.local_init_done
		.local_cal_success          (mem_if_ddr3_emif_0_status_local_cal_success),                   //                   .local_cal_success
		.local_cal_fail             (mem_if_ddr3_emif_0_status_local_cal_fail),                      //                   .local_cal_fail
		.oct_rzqin                  (oct_rzqin),                                                     //                oct.rzqin
		.pll_mem_clk                (),                                                              //        pll_sharing.pll_mem_clk
		.pll_write_clk              (),                                                              //                   .pll_write_clk
		.pll_locked                 (),                                                              //                   .pll_locked
		.pll_write_clk_pre_phy_clk  (),                                                              //                   .pll_write_clk_pre_phy_clk
		.pll_addr_cmd_clk           (),                                                              //                   .pll_addr_cmd_clk
		.pll_avl_clk                (),                                                              //                   .pll_avl_clk
		.pll_config_clk             (),                                                              //                   .pll_config_clk
		.pll_mem_phy_clk            (),                                                              //                   .pll_mem_phy_clk
		.afi_phy_clk                (),                                                              //                   .afi_phy_clk
		.pll_avl_phy_clk            ()                                                               //                   .pll_avl_phy_clk
	);

	top_mipi_pwdn_n mipi_pwdn_n (
		.clk        (pll_0_outclk0_clk),                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_1_mipi_pwdn_n_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_mipi_pwdn_n_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_mipi_pwdn_n_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_mipi_pwdn_n_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_mipi_pwdn_n_s1_readdata),   //                    .readdata
		.out_port   (mipi_pwdn_n_external_connection_export)       // external_connection.export
	);

	top_mipi_pwdn_n mipi_reset_n (
		.clk        (pll_0_outclk0_clk),                            //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_1_mipi_reset_n_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_mipi_reset_n_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_mipi_reset_n_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_mipi_reset_n_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_mipi_reset_n_s1_readdata),   //                    .readdata
		.out_port   (mipi_reset_n_external_connection_export)       // external_connection.export
	);

	top_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (pll_0_outclk0_clk),                                          //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                            //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nios2_gen2_0_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_gen2_0_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                           //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	top_nios_ram nios_ram (
		.clk        (pll_0_outclk0_clk),                        //   clk1.clk
		.address    (mm_interconnect_1_nios_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_1_nios_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_1_nios_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_1_nios_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_1_nios_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_1_nios_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_1_nios_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),           // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),       //       .reset_req
		.freeze     (1'b0)                                      // (terminated)
	);

	top_ocm_256k_dma ocm_256k_dma (
		.clk         (pll_0_outclk0_clk),                            //   clk1.clk
		.address     (mm_interconnect_1_ocm_256k_dma_s1_address),    //     s1.address
		.clken       (mm_interconnect_1_ocm_256k_dma_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_1_ocm_256k_dma_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_1_ocm_256k_dma_s1_write),      //       .write
		.readdata    (mm_interconnect_1_ocm_256k_dma_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_1_ocm_256k_dma_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_1_ocm_256k_dma_s1_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),               // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),           //       .reset_req
		.address2    (mm_interconnect_2_ocm_256k_dma_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_2_ocm_256k_dma_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_2_ocm_256k_dma_s2_clken),      //       .clken
		.write2      (mm_interconnect_2_ocm_256k_dma_s2_write),      //       .write
		.readdata2   (mm_interconnect_2_ocm_256k_dma_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_2_ocm_256k_dma_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_2_ocm_256k_dma_s2_byteenable), //       .byteenable
		.clk2        (pcie_256_dma_coreclkout_clk),                  //   clk2.clk
		.reset2      (rst_controller_002_reset_out_reset),           // reset2.reset
		.reset_req2  (rst_controller_002_reset_out_reset_req),       //       .reset_req
		.freeze      (1'b0)                                          // (terminated)
	);

	altpcie_256_hip_avmm_hwtcl #(
		.INTENDED_DEVICE_FAMILY                   ("Cyclone V"),
		.lane_mask_hwtcl                          ("x4"),
		.gen123_lane_rate_mode_hwtcl              ("Gen2 (5.0 Gbps)"),
		.DMA_WIDTH                                (128),
		.DMA_BE_WIDTH                             (16),
		.DMA_BRST_CNT_W                           (6),
		.port_type_hwtcl                          ("Native endpoint"),
		.pcie_spec_version_hwtcl                  ("2.1"),
		.pll_refclk_freq_hwtcl                    ("100 MHz"),
		.set_pld_clk_x1_625MHz_hwtcl              (0),
		.internal_controller_hwtcl                (1),
		.enable_cra_hwtcl                         (0),
		.enable_rxm_burst_hwtcl                   (0),
		.in_cvp_mode_hwtcl                        (0),
		.enable_tl_only_sim_hwtcl                 (0),
		.use_atx_pll_hwtcl                        (0),
		.dma_use_scfifo_ext_hwtcl                 (0),
		.bar0_type_hwtcl                          (64),
		.bar0_size_mask_hwtcl                     (9),
		.bar0_io_space_hwtcl                      ("Disabled"),
		.bar0_64bit_mem_space_hwtcl               ("Enabled"),
		.bar0_prefetchable_hwtcl                  ("Enabled"),
		.bar1_type_hwtcl                          (1),
		.bar1_size_mask_hwtcl                     (0),
		.bar1_io_space_hwtcl                      ("Disabled"),
		.bar1_prefetchable_hwtcl                  ("Disabled"),
		.bar2_type_hwtcl                          (64),
		.bar2_size_mask_hwtcl                     (31),
		.bar2_io_space_hwtcl                      ("Disabled"),
		.bar2_64bit_mem_space_hwtcl               ("Enabled"),
		.bar2_prefetchable_hwtcl                  ("Enabled"),
		.bar3_type_hwtcl                          (1),
		.bar3_size_mask_hwtcl                     (0),
		.bar3_io_space_hwtcl                      ("Disabled"),
		.bar3_prefetchable_hwtcl                  ("Disabled"),
		.bar4_type_hwtcl                          (1),
		.bar4_size_mask_hwtcl                     (0),
		.bar4_io_space_hwtcl                      ("Disabled"),
		.bar4_64bit_mem_space_hwtcl               ("Disabled"),
		.bar4_prefetchable_hwtcl                  ("Disabled"),
		.bar5_type_hwtcl                          (1),
		.bar5_size_mask_hwtcl                     (0),
		.rd_dma_size_mask_hwtcl                   (32),
		.wr_dma_size_mask_hwtcl                   (31),
		.bar5_io_space_hwtcl                      ("Disabled"),
		.bar5_prefetchable_hwtcl                  ("Disabled"),
		.vendor_id_hwtcl                          (4466),
		.device_id_hwtcl                          (57347),
		.revision_id_hwtcl                        (1),
		.class_code_hwtcl                         (0),
		.subsystem_vendor_id_hwtcl                (4369),
		.subsystem_device_id_hwtcl                (13409),
		.max_payload_size_hwtcl                   (256),
		.extend_tag_field_hwtcl                   ("32"),
		.completion_timeout_hwtcl                 ("ABCD"),
		.enable_completion_timeout_disable_hwtcl  (1),
		.use_aer_hwtcl                            (0),
		.ecrc_check_capable_hwtcl                 (0),
		.ecrc_gen_capable_hwtcl                   (0),
		.use_crc_forwarding_hwtcl                 (0),
		.port_link_number_hwtcl                   (1),
		.dll_active_report_support_hwtcl          (0),
		.surprise_down_error_support_hwtcl        (0),
		.slotclkcfg_hwtcl                         (1),
		.msi_multi_message_capable_hwtcl          ("1"),
		.msi_64bit_addressing_capable_hwtcl       ("true"),
		.msi_masking_capable_hwtcl                ("false"),
		.msi_support_hwtcl                        ("true"),
		.enable_function_msix_support_hwtcl       (0),
		.msix_table_size_hwtcl                    (0),
		.msix_table_offset_hwtcl                  ("0"),
		.msix_table_bir_hwtcl                     (0),
		.msix_pba_offset_hwtcl                    ("0"),
		.msix_pba_bir_hwtcl                       (0),
		.enable_slot_register_hwtcl               (0),
		.slot_power_scale_hwtcl                   (0),
		.slot_power_limit_hwtcl                   (0),
		.slot_number_hwtcl                        (0),
		.endpoint_l0_latency_hwtcl                (0),
		.endpoint_l1_latency_hwtcl                (0),
		.avmm_width_hwtcl                         (256),
		.avmm_burst_width_hwtcl                   (7),
		.TX_S_ADDR_WIDTH                          (64),
		.ast_width_hwtcl                          ("Avalon-ST 128-bit"),
		.use_ast_parity                           (0),
		.millisecond_cycle_count_hwtcl            (124250),
		.set_pll_coreclkout_cout_hwtcl            ("NA"),
		.set_pll_coreclkout_cin_hwtcl             ("NA"),
		.port_width_be_hwtcl                      (16),
		.port_width_data_hwtcl                    (128),
		.hip_reconfig_hwtcl                       (0),
		.vsec_id_hwtcl                            (40960),
		.vsec_rev_hwtcl                           (0),
		.expansion_base_address_register_hwtcl    (0),
		.prefetchable_mem_window_addr_width_hwtcl (0),
		.bypass_cdc_hwtcl                         ("false"),
		.enable_rx_buffer_checking_hwtcl          ("false"),
		.disable_link_x2_support_hwtcl            ("false"),
		.wrong_device_id_hwtcl                    ("disable"),
		.data_pack_rx_hwtcl                       ("disable"),
		.ltssm_1ms_timeout_hwtcl                  ("disable"),
		.ltssm_freqlocked_check_hwtcl             ("disable"),
		.deskew_comma_hwtcl                       ("skp_eieos_deskw"),
		.device_number_hwtcl                      (0),
		.pipex1_debug_sel_hwtcl                   ("disable"),
		.pclk_out_sel_hwtcl                       ("pclk"),
		.no_soft_reset_hwtcl                      ("false"),
		.maximum_current_hwtcl                    (0),
		.d1_support_hwtcl                         ("false"),
		.d2_support_hwtcl                         ("false"),
		.d0_pme_hwtcl                             ("false"),
		.d1_pme_hwtcl                             ("false"),
		.d2_pme_hwtcl                             ("false"),
		.d3_hot_pme_hwtcl                         ("false"),
		.d3_cold_pme_hwtcl                        ("false"),
		.low_priority_vc_hwtcl                    ("single_vc"),
		.disable_snoop_packet_hwtcl               ("false"),
		.enable_l1_aspm_hwtcl                     ("false"),
		.rx_ei_l0s_hwtcl                          (0),
		.enable_l0s_aspm_hwtcl                    ("false"),
		.aspm_config_management_hwtcl             ("true"),
		.l1_exit_latency_sameclock_hwtcl          (0),
		.l1_exit_latency_diffclock_hwtcl          (0),
		.hot_plug_support_hwtcl                   (0),
		.extended_tag_reset_hwtcl                 ("false"),
		.no_command_completed_hwtcl               ("false"),
		.interrupt_pin_hwtcl                      ("inta"),
		.bridge_port_vga_enable_hwtcl             ("false"),
		.bridge_port_ssid_support_hwtcl           ("false"),
		.ssvid_hwtcl                              (0),
		.ssid_hwtcl                               (0),
		.eie_before_nfts_count_hwtcl              (4),
		.gen2_diffclock_nfts_count_hwtcl          (255),
		.gen2_sameclock_nfts_count_hwtcl          (255),
		.l0_exit_latency_sameclock_hwtcl          (6),
		.l0_exit_latency_diffclock_hwtcl          (6),
		.atomic_op_routing_hwtcl                  ("false"),
		.atomic_op_completer_32bit_hwtcl          ("false"),
		.atomic_op_completer_64bit_hwtcl          ("false"),
		.cas_completer_128bit_hwtcl               ("false"),
		.ltr_mechanism_hwtcl                      ("false"),
		.tph_completer_hwtcl                      ("false"),
		.extended_format_field_hwtcl              ("false"),
		.atomic_malformed_hwtcl                   ("true"),
		.flr_capability_hwtcl                     ("false"),
		.enable_adapter_half_rate_mode_hwtcl      ("true"),
		.vc0_clk_enable_hwtcl                     ("true"),
		.register_pipe_signals_hwtcl              ("true"),
		.skp_os_gen3_count_hwtcl                  (0),
		.tx_cdc_almost_empty_hwtcl                (5),
		.rx_l0s_count_idl_hwtcl                   (0),
		.cdc_dummy_insert_limit_hwtcl             (11),
		.ei_delay_powerdown_count_hwtcl           (10),
		.skp_os_schedule_count_hwtcl              (0),
		.fc_init_timer_hwtcl                      (1024),
		.l01_entry_latency_hwtcl                  (31),
		.flow_control_update_count_hwtcl          (30),
		.flow_control_timeout_count_hwtcl         (200),
		.retry_buffer_last_active_address_hwtcl   (2047),
		.reserved_debug_hwtcl                     (0),
		.bypass_clk_switch_hwtcl                  ("disable"),
		.l2_async_logic_hwtcl                     ("disable"),
		.indicator_hwtcl                          (0),
		.diffclock_nfts_count_hwtcl               (128),
		.sameclock_nfts_count_hwtcl               (128),
		.rx_cdc_almost_full_hwtcl                 (12),
		.tx_cdc_almost_full_hwtcl                 (11),
		.credit_buffer_allocation_aux_hwtcl       ("balanced"),
		.vc0_rx_flow_ctrl_posted_header_hwtcl     (16),
		.vc0_rx_flow_ctrl_posted_data_hwtcl       (16),
		.vc0_rx_flow_ctrl_nonposted_header_hwtcl  (16),
		.vc0_rx_flow_ctrl_nonposted_data_hwtcl    (0),
		.vc0_rx_flow_ctrl_compl_header_hwtcl      (0),
		.vc0_rx_flow_ctrl_compl_data_hwtcl        (0),
		.cpl_spc_header_hwtcl                     (67),
		.cpl_spc_data_hwtcl                       (269),
		.gen3_rxfreqlock_counter_hwtcl            (0),
		.gen3_skip_ph2_ph3_hwtcl                  (0),
		.g3_bypass_equlz_hwtcl                    (0),
		.cvp_data_compressed_hwtcl                ("false"),
		.cvp_data_encrypted_hwtcl                 ("false"),
		.cvp_mode_reset_hwtcl                     ("false"),
		.cvp_clk_reset_hwtcl                      ("false"),
		.cseb_cpl_status_during_cvp_hwtcl         ("config_retry_status"),
		.core_clk_sel_hwtcl                       ("pld_clk"),
		.cvp_rate_sel_hwtcl                       ("full_rate"),
		.g3_dis_rx_use_prst_hwtcl                 ("true"),
		.g3_dis_rx_use_prst_ep_hwtcl              ("true"),
		.deemphasis_enable_hwtcl                  ("false"),
		.reconfig_to_xcvr_width                   (350),
		.reconfig_from_xcvr_width                 (230),
		.single_rx_detect_hwtcl                   (4),
		.hip_hard_reset_hwtcl                     (1),
		.use_cvp_update_core_pof_hwtcl            (0),
		.pcie_inspector_hwtcl                     (0),
		.tlp_inspector_hwtcl                      (0),
		.tlp_inspector_use_signal_probe_hwtcl     (0),
		.tlp_insp_trg_dw0_hwtcl                   (2049),
		.tlp_insp_trg_dw1_hwtcl                   (0),
		.tlp_insp_trg_dw2_hwtcl                   (0),
		.tlp_insp_trg_dw3_hwtcl                   (0),
		.use_tl_cfg_sync_hwtcl                    (1),
		.hwtcl_override_g2_txvod                  (1),
		.rpre_emph_a_val_hwtcl                    (9),
		.rpre_emph_b_val_hwtcl                    (0),
		.rpre_emph_c_val_hwtcl                    (16),
		.rpre_emph_d_val_hwtcl                    (13),
		.rpre_emph_e_val_hwtcl                    (5),
		.rvod_sel_a_val_hwtcl                     (42),
		.rvod_sel_b_val_hwtcl                     (38),
		.rvod_sel_c_val_hwtcl                     (38),
		.rvod_sel_d_val_hwtcl                     (43),
		.rvod_sel_e_val_hwtcl                     (15),
		.av_rpre_emph_a_val_hwtcl                 (12),
		.av_rpre_emph_b_val_hwtcl                 (0),
		.av_rpre_emph_c_val_hwtcl                 (19),
		.av_rpre_emph_d_val_hwtcl                 (13),
		.av_rpre_emph_e_val_hwtcl                 (21),
		.av_rvod_sel_a_val_hwtcl                  (42),
		.av_rvod_sel_b_val_hwtcl                  (30),
		.av_rvod_sel_c_val_hwtcl                  (43),
		.av_rvod_sel_d_val_hwtcl                  (43),
		.av_rvod_sel_e_val_hwtcl                  (9),
		.cv_rpre_emph_a_val_hwtcl                 (11),
		.cv_rpre_emph_b_val_hwtcl                 (0),
		.cv_rpre_emph_c_val_hwtcl                 (22),
		.cv_rpre_emph_d_val_hwtcl                 (12),
		.cv_rpre_emph_e_val_hwtcl                 (21),
		.cv_rvod_sel_a_val_hwtcl                  (50),
		.cv_rvod_sel_b_val_hwtcl                  (34),
		.cv_rvod_sel_c_val_hwtcl                  (50),
		.cv_rvod_sel_d_val_hwtcl                  (50),
		.cv_rvod_sel_e_val_hwtcl                  (9)
	) pcie_256_dma (
		.coreclkout           (pcie_256_dma_coreclkout_clk),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //          coreclkout.clk
		.refclk               (refclk_clk),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //              refclk.clk
		.npor                 (pcie_rstn_npor),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //                npor.npor
		.pin_perst            (pcie_rstn_pin_perst),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                    .pin_perst
		.reset_status         (pcie_256_dma_nreset_status_reset),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //       nreset_status.reset_n
		.RxmAddress_2_o       (pcie_256_dma_rxm_bar2_address),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //            Rxm_BAR2.address
		.RxmRead_2_o          (pcie_256_dma_rxm_bar2_read),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //                    .read
		.RxmWaitRequest_2_i   (pcie_256_dma_rxm_bar2_waitrequest),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .waitrequest
		.RxmWrite_2_o         (pcie_256_dma_rxm_bar2_write),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                    .write
		.RxmReadDataValid_2_i (pcie_256_dma_rxm_bar2_readdatavalid),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                    .readdatavalid
		.RxmReadData_2_i      (pcie_256_dma_rxm_bar2_readdata),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //                    .readdata
		.RxmWriteData_2_o     (pcie_256_dma_rxm_bar2_writedata),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //                    .writedata
		.RxmByteEnable_2_o    (pcie_256_dma_rxm_bar2_byteenable),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .byteenable
		.TxsAddress_i         (mm_interconnect_4_pcie_256_dma_txs_address),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //                 Txs.address
		.TxsChipSelect_i      (mm_interconnect_4_pcie_256_dma_txs_chipselect),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //                    .chipselect
		.TxsByteEnable_i      (mm_interconnect_4_pcie_256_dma_txs_byteenable),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //                    .byteenable
		.TxsReadData_o        (mm_interconnect_4_pcie_256_dma_txs_readdata),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                    .readdata
		.TxsWriteData_i       (mm_interconnect_4_pcie_256_dma_txs_writedata),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //                    .writedata
		.TxsRead_i            (mm_interconnect_4_pcie_256_dma_txs_read),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                    .read
		.TxsWrite_i           (mm_interconnect_4_pcie_256_dma_txs_write),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                    .write
		.TxsReadDataValid_o   (mm_interconnect_4_pcie_256_dma_txs_readdatavalid),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .readdatavalid
		.TxsWaitRequest_o     (mm_interconnect_4_pcie_256_dma_txs_waitrequest),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //                    .waitrequest
		.RdDmaAddress_o       (pcie_256_dma_dma_rd_master_address),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //       dma_rd_master.address
		.RdDmaWrite_o         (pcie_256_dma_dma_rd_master_write),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .write
		.RdDmaWriteData_o     (pcie_256_dma_dma_rd_master_writedata),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .writedata
		.RdDmaWaitRequest_i   (pcie_256_dma_dma_rd_master_waitrequest),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //                    .waitrequest
		.RdDmaBurstCount_o    (pcie_256_dma_dma_rd_master_burstcount),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //                    .burstcount
		.RdDmaWriteEnable_o   (pcie_256_dma_dma_rd_master_byteenable),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //                    .byteenable
		.WrDmaAddress_o       (pcie_256_dma_dma_wr_master_address),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //       dma_wr_master.address
		.WrDmaRead_o          (pcie_256_dma_dma_wr_master_read),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //                    .read
		.WrDmaWaitRequest_i   (pcie_256_dma_dma_wr_master_waitrequest),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //                    .waitrequest
		.WrDmaBurstCount_o    (pcie_256_dma_dma_wr_master_burstcount),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //                    .burstcount
		.WrDmaReadDataValid_i (pcie_256_dma_dma_wr_master_readdatavalid),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                    .readdatavalid
		.WrDmaReadData_i      (pcie_256_dma_dma_wr_master_readdata),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                    .readdata
		.WrDTSChipSelect_i    (mm_interconnect_2_pcie_256_dma_wr_dts_slave_chipselect),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //        wr_dts_slave.chipselect
		.WrDTSWrite_i         (mm_interconnect_2_pcie_256_dma_wr_dts_slave_write),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .write
		.WrDTSBurstCount_i    (mm_interconnect_2_pcie_256_dma_wr_dts_slave_burstcount),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //                    .burstcount
		.WrDTSAddress_i       (mm_interconnect_2_pcie_256_dma_wr_dts_slave_address),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                    .address
		.WrDTSWriteData_i     (mm_interconnect_2_pcie_256_dma_wr_dts_slave_writedata),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //                    .writedata
		.WrDTSWaitRequest_o   (mm_interconnect_2_pcie_256_dma_wr_dts_slave_waitrequest),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                    .waitrequest
		.RdDTSChipSelect_i    (mm_interconnect_2_pcie_256_dma_rd_dts_slave_chipselect),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //        rd_dts_slave.chipselect
		.RdDTSWrite_i         (mm_interconnect_2_pcie_256_dma_rd_dts_slave_write),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .write
		.RdDTSBurstCount_i    (mm_interconnect_2_pcie_256_dma_rd_dts_slave_burstcount),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //                    .burstcount
		.RdDTSAddress_i       (mm_interconnect_2_pcie_256_dma_rd_dts_slave_address),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                    .address
		.RdDTSWriteData_i     (mm_interconnect_2_pcie_256_dma_rd_dts_slave_writedata),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //                    .writedata
		.RdDTSWaitRequest_o   (mm_interconnect_2_pcie_256_dma_rd_dts_slave_waitrequest),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                    .waitrequest
		.WrDCMAddress_o       (pcie_256_dma_wr_dcm_master_address),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //       wr_dcm_master.address
		.WrDCMWrite_o         (pcie_256_dma_wr_dcm_master_write),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .write
		.WrDCMWriteData_o     (pcie_256_dma_wr_dcm_master_writedata),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .writedata
		.WrDCMRead_o          (pcie_256_dma_wr_dcm_master_read),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //                    .read
		.WrDCMByteEnable_o    (pcie_256_dma_wr_dcm_master_byteenable),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //                    .byteenable
		.WrDCMWaitRequest_i   (pcie_256_dma_wr_dcm_master_waitrequest),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //                    .waitrequest
		.WrDCMReadData_i      (pcie_256_dma_wr_dcm_master_readdata),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                    .readdata
		.WrDCMReadDataValid_i (pcie_256_dma_wr_dcm_master_readdatavalid),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                    .readdatavalid
		.RdDCMAddress_o       (pcie_256_dma_rd_dcm_master_address),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //       rd_dcm_master.address
		.RdDCMWrite_o         (pcie_256_dma_rd_dcm_master_write),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .write
		.RdDCMWriteData_o     (pcie_256_dma_rd_dcm_master_writedata),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .writedata
		.RdDCMRead_o          (pcie_256_dma_rd_dcm_master_read),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //                    .read
		.RdDCMByteEnable_o    (pcie_256_dma_rd_dcm_master_byteenable),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //                    .byteenable
		.RdDCMWaitRequest_i   (pcie_256_dma_rd_dcm_master_waitrequest),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //                    .waitrequest
		.RdDCMReadData_i      (pcie_256_dma_rd_dcm_master_readdata),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                    .readdata
		.RdDCMReadDataValid_i (pcie_256_dma_rd_dcm_master_readdatavalid),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                    .readdatavalid
		.IntxReq_i            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //      INTX_Interface.intx_req
		.IntxAck_o            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .intx_ack
		.MsiIntfc_o           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //       MSI_Interface.msi_intfc
		.MsixIntfc_o          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //      MSIX_Interface.msix_intfc
		.reconfig_to_xcvr     (alt_xcvr_reconfig_0_reconfig_to_xcvr_reconfig_to_xcvr),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //    reconfig_to_xcvr.reconfig_to_xcvr
		.reconfig_from_xcvr   (pcie_256_dma_reconfig_from_xcvr_reconfig_from_xcvr),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //  reconfig_from_xcvr.reconfig_from_xcvr
		.fixedclk_locked      (pcie_256_hip_avmm_0_reconfig_clk_locked_fixedclk_locked),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         // reconfig_clk_locked.fixedclk_locked
		.rx_in0               (hip_serial_rx_in0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //          hip_serial.rx_in0
		.rx_in1               (hip_serial_rx_in1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .rx_in1
		.rx_in2               (hip_serial_rx_in2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .rx_in2
		.rx_in3               (hip_serial_rx_in3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .rx_in3
		.tx_out0              (hip_serial_tx_out0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                    .tx_out0
		.tx_out1              (hip_serial_tx_out1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                    .tx_out1
		.tx_out2              (hip_serial_tx_out2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                    .tx_out2
		.tx_out3              (hip_serial_tx_out3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                    .tx_out3
		.sim_pipe_pclk_in     (hip_pipe_sim_pipe_pclk_in),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //            hip_pipe.sim_pipe_pclk_in
		.sim_pipe_rate        (hip_pipe_sim_pipe_rate),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //                    .sim_pipe_rate
		.sim_ltssmstate       (hip_pipe_sim_ltssmstate),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                    .sim_ltssmstate
		.eidleinfersel0       (hip_pipe_eidleinfersel0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                    .eidleinfersel0
		.eidleinfersel1       (hip_pipe_eidleinfersel1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                    .eidleinfersel1
		.eidleinfersel2       (hip_pipe_eidleinfersel2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                    .eidleinfersel2
		.eidleinfersel3       (hip_pipe_eidleinfersel3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                    .eidleinfersel3
		.powerdown0           (hip_pipe_powerdown0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                    .powerdown0
		.powerdown1           (hip_pipe_powerdown1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                    .powerdown1
		.powerdown2           (hip_pipe_powerdown2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                    .powerdown2
		.powerdown3           (hip_pipe_powerdown3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                    .powerdown3
		.rxpolarity0          (hip_pipe_rxpolarity0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .rxpolarity0
		.rxpolarity1          (hip_pipe_rxpolarity1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .rxpolarity1
		.rxpolarity2          (hip_pipe_rxpolarity2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .rxpolarity2
		.rxpolarity3          (hip_pipe_rxpolarity3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .rxpolarity3
		.txcompl0             (hip_pipe_txcompl0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .txcompl0
		.txcompl1             (hip_pipe_txcompl1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .txcompl1
		.txcompl2             (hip_pipe_txcompl2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .txcompl2
		.txcompl3             (hip_pipe_txcompl3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .txcompl3
		.txdata0              (hip_pipe_txdata0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .txdata0
		.txdata1              (hip_pipe_txdata1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .txdata1
		.txdata2              (hip_pipe_txdata2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .txdata2
		.txdata3              (hip_pipe_txdata3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .txdata3
		.txdatak0             (hip_pipe_txdatak0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .txdatak0
		.txdatak1             (hip_pipe_txdatak1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .txdatak1
		.txdatak2             (hip_pipe_txdatak2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .txdatak2
		.txdatak3             (hip_pipe_txdatak3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .txdatak3
		.txdetectrx0          (hip_pipe_txdetectrx0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .txdetectrx0
		.txdetectrx1          (hip_pipe_txdetectrx1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .txdetectrx1
		.txdetectrx2          (hip_pipe_txdetectrx2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .txdetectrx2
		.txdetectrx3          (hip_pipe_txdetectrx3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .txdetectrx3
		.txelecidle0          (hip_pipe_txelecidle0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .txelecidle0
		.txelecidle1          (hip_pipe_txelecidle1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .txelecidle1
		.txelecidle2          (hip_pipe_txelecidle2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .txelecidle2
		.txelecidle3          (hip_pipe_txelecidle3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .txelecidle3
		.txdeemph0            (hip_pipe_txdeemph0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                    .txdeemph0
		.txdeemph1            (hip_pipe_txdeemph1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                    .txdeemph1
		.txdeemph2            (hip_pipe_txdeemph2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                    .txdeemph2
		.txdeemph3            (hip_pipe_txdeemph3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                    .txdeemph3
		.txmargin0            (hip_pipe_txmargin0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                    .txmargin0
		.txmargin1            (hip_pipe_txmargin1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                    .txmargin1
		.txmargin2            (hip_pipe_txmargin2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                    .txmargin2
		.txmargin3            (hip_pipe_txmargin3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                    .txmargin3
		.txswing0             (hip_pipe_txswing0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .txswing0
		.txswing1             (hip_pipe_txswing1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .txswing1
		.txswing2             (hip_pipe_txswing2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .txswing2
		.txswing3             (hip_pipe_txswing3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .txswing3
		.phystatus0           (hip_pipe_phystatus0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                    .phystatus0
		.phystatus1           (hip_pipe_phystatus1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                    .phystatus1
		.phystatus2           (hip_pipe_phystatus2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                    .phystatus2
		.phystatus3           (hip_pipe_phystatus3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                    .phystatus3
		.rxdata0              (hip_pipe_rxdata0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .rxdata0
		.rxdata1              (hip_pipe_rxdata1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .rxdata1
		.rxdata2              (hip_pipe_rxdata2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .rxdata2
		.rxdata3              (hip_pipe_rxdata3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .rxdata3
		.rxdatak0             (hip_pipe_rxdatak0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .rxdatak0
		.rxdatak1             (hip_pipe_rxdatak1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .rxdatak1
		.rxdatak2             (hip_pipe_rxdatak2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .rxdatak2
		.rxdatak3             (hip_pipe_rxdatak3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .rxdatak3
		.rxelecidle0          (hip_pipe_rxelecidle0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .rxelecidle0
		.rxelecidle1          (hip_pipe_rxelecidle1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .rxelecidle1
		.rxelecidle2          (hip_pipe_rxelecidle2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .rxelecidle2
		.rxelecidle3          (hip_pipe_rxelecidle3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                    .rxelecidle3
		.rxstatus0            (hip_pipe_rxstatus0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                    .rxstatus0
		.rxstatus1            (hip_pipe_rxstatus1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                    .rxstatus1
		.rxstatus2            (hip_pipe_rxstatus2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                    .rxstatus2
		.rxstatus3            (hip_pipe_rxstatus3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                    .rxstatus3
		.rxvalid0             (hip_pipe_rxvalid0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .rxvalid0
		.rxvalid1             (hip_pipe_rxvalid1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .rxvalid1
		.rxvalid2             (hip_pipe_rxvalid2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .rxvalid2
		.rxvalid3             (hip_pipe_rxvalid3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                    .rxvalid3
		.test_in              (hip_ctrl_test_in),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //            hip_ctrl.test_in
		.simu_mode_pipe       (hip_ctrl_simu_mode_pipe),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                    .simu_mode_pipe
		.derr_cor_ext_rcv     (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //          hip_status.derr_cor_ext_rcv
		.derr_cor_ext_rpl     (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .derr_cor_ext_rpl
		.derr_rpl             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .derr_rpl
		.dlup_exit            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .dlup_exit
		.ev128ns              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .ev128ns
		.ev1us                (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .ev1us
		.hotrst_exit          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .hotrst_exit
		.int_status           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .int_status
		.l2_exit              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .l2_exit
		.lane_act             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .lane_act
		.ltssmstate           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .ltssmstate
		.ko_cpl_spc_header    (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .ko_cpl_spc_header
		.ko_cpl_spc_data      (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .ko_cpl_spc_data
		.currentspeed         (pcie_256_dma_hip_currentspeed_currentspeed),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //    hip_currentspeed.currentspeed
		.tl_cfg_add           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //           config_tl.tl_cfg_add
		.tl_cfg_ctl           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .tl_cfg_ctl
		.tl_cfg_sts           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                    .tl_cfg_sts
		.RdDmaRxValid_i       (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.RdDmaRxData_i        (160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //         (terminated)
		.RdDmaRxReady_o       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.RdDmaTxData_o        (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.RdDmaTxValid_o       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.WrDmaRxValid_i       (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.WrDmaRxData_i        (160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //         (terminated)
		.WrDmaRxReady_o       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.WrDmaTxData_o        (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.WrDmaTxValid_o       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.rx_in4               (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rx_in5               (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rx_in6               (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rx_in7               (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.tx_out4              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.tx_out5              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.tx_out6              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.tx_out7              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.eidleinfersel4       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.eidleinfersel5       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.eidleinfersel6       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.eidleinfersel7       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.powerdown4           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.powerdown5           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.powerdown6           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.powerdown7           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.rxpolarity4          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.rxpolarity5          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.rxpolarity6          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.rxpolarity7          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txcompl4             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txcompl5             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txcompl6             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txcompl7             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txdata4              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txdata5              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txdata6              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txdata7              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txdatak4             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txdatak5             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txdatak6             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txdatak7             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txdetectrx4          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txdetectrx5          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txdetectrx6          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txdetectrx7          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txelecidle4          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txelecidle5          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txelecidle6          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txelecidle7          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txdeemph4            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txdeemph5            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txdeemph6            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txdeemph7            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txmargin4            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txmargin5            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txmargin6            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txmargin7            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txswing4             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txswing5             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txswing6             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txswing7             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.phystatus4           (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.phystatus5           (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.phystatus6           (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.phystatus7           (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxdata4              (8'b00000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //         (terminated)
		.rxdata5              (8'b00000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //         (terminated)
		.rxdata6              (8'b00000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //         (terminated)
		.rxdata7              (8'b00000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //         (terminated)
		.rxdatak4             (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxdatak5             (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxdatak6             (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxdatak7             (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxelecidle4          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxelecidle5          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxelecidle6          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxelecidle7          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxstatus4            (3'b000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //         (terminated)
		.rxstatus5            (3'b000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //         (terminated)
		.rxstatus6            (3'b000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //         (terminated)
		.rxstatus7            (3'b000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //         (terminated)
		.rxvalid4             (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxvalid5             (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxvalid6             (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxvalid7             (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxdataskip0          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxdataskip1          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxdataskip2          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxdataskip3          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxdataskip4          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxdataskip5          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxdataskip6          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxdataskip7          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxblkst0             (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxblkst1             (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxblkst2             (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxblkst3             (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxblkst4             (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxblkst5             (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxblkst6             (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxblkst7             (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxsynchd0            (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //         (terminated)
		.rxsynchd1            (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //         (terminated)
		.rxsynchd2            (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //         (terminated)
		.rxsynchd3            (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //         (terminated)
		.rxsynchd4            (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //         (terminated)
		.rxsynchd5            (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //         (terminated)
		.rxsynchd6            (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //         (terminated)
		.rxsynchd7            (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //         (terminated)
		.rxfreqlocked0        (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxfreqlocked1        (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxfreqlocked2        (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxfreqlocked3        (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxfreqlocked4        (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxfreqlocked5        (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxfreqlocked6        (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.rxfreqlocked7        (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //         (terminated)
		.currentcoeff0        (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.currentcoeff1        (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.currentcoeff2        (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.currentcoeff3        (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.currentcoeff4        (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.currentcoeff5        (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.currentcoeff6        (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.currentcoeff7        (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.currentrxpreset0     (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.currentrxpreset1     (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.currentrxpreset2     (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.currentrxpreset3     (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.currentrxpreset4     (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.currentrxpreset5     (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.currentrxpreset6     (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.currentrxpreset7     (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txsynchd0            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txsynchd1            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txsynchd2            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txsynchd3            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txsynchd4            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txsynchd5            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txsynchd6            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txsynchd7            (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txblkst0             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txblkst1             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txblkst2             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txblkst3             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txblkst4             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txblkst5             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txblkst6             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.txblkst7             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.tlbfm_in             (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.tlbfm_out            (1001'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000), //         (terminated)
		.dlup                 (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.rx_par_err           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.tx_par_err           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         (terminated)
		.cfg_par_err          ()                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //         (terminated)
	);

	altpcie_reconfig_driver #(
		.INTENDED_DEVICE_FAMILY        ("Cyclone V"),
		.gen123_lane_rate_mode_hwtcl   ("Gen2 (5.0 Gbps)"),
		.number_of_reconfig_interfaces (5)
	) pcie_reconfig_driver_0 (
		.reconfig_xcvr_clk         (pcie_256_dma_coreclkout_clk),                      // reconfig_xcvr_clk.clk
		.reconfig_xcvr_rst         (rst_controller_002_reset_out_reset),               // reconfig_xcvr_rst.reset
		.reconfig_mgmt_address     (pcie_reconfig_driver_0_reconfig_mgmt_address),     //     reconfig_mgmt.address
		.reconfig_mgmt_read        (pcie_reconfig_driver_0_reconfig_mgmt_read),        //                  .read
		.reconfig_mgmt_readdata    (pcie_reconfig_driver_0_reconfig_mgmt_readdata),    //                  .readdata
		.reconfig_mgmt_waitrequest (pcie_reconfig_driver_0_reconfig_mgmt_waitrequest), //                  .waitrequest
		.reconfig_mgmt_write       (pcie_reconfig_driver_0_reconfig_mgmt_write),       //                  .write
		.reconfig_mgmt_writedata   (pcie_reconfig_driver_0_reconfig_mgmt_writedata),   //                  .writedata
		.currentspeed              (pcie_256_dma_hip_currentspeed_currentspeed),       //  hip_currentspeed.currentspeed
		.reconfig_busy             (),                                                 //     reconfig_busy.reconfig_busy
		.pld_clk                   (pcie_256_dma_coreclkout_clk),                      //           pld_clk.clk
		.derr_cor_ext_rcv_drv      (),                                                 //    hip_status_drv.derr_cor_ext_rcv
		.derr_cor_ext_rpl_drv      (),                                                 //                  .derr_cor_ext_rpl
		.derr_rpl_drv              (),                                                 //                  .derr_rpl
		.dlup_exit_drv             (),                                                 //                  .dlup_exit
		.ev128ns_drv               (),                                                 //                  .ev128ns
		.ev1us_drv                 (),                                                 //                  .ev1us
		.hotrst_exit_drv           (),                                                 //                  .hotrst_exit
		.int_status_drv            (),                                                 //                  .int_status
		.l2_exit_drv               (),                                                 //                  .l2_exit
		.lane_act_drv              (),                                                 //                  .lane_act
		.ltssmstate_drv            (),                                                 //                  .ltssmstate
		.ko_cpl_spc_header_drv     (),                                                 //                  .ko_cpl_spc_header
		.ko_cpl_spc_data_drv       (),                                                 //                  .ko_cpl_spc_data
		.cal_busy_in               (),                                                 //       (terminated)
		.dlup_drv                  (1'b0),                                             //       (terminated)
		.rx_par_err_drv            (1'b0),                                             //       (terminated)
		.tx_par_err_drv            (2'b00),                                            //       (terminated)
		.cfg_par_err_drv           (1'b0)                                              //       (terminated)
	);

	top_pio_button pio_button (
		.clk        (pll_0_outclk0_clk),                          //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_1_pio_button_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_pio_button_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_pio_button_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_pio_button_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_pio_button_s1_readdata),   //                    .readdata
		.in_port    (pio_button_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver4_irq)                    //                 irq.irq
	);

	top_pio_led pio_led (
		.clk        (pll_0_outclk0_clk),                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_1_pio_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_pio_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_pio_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_pio_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_pio_led_s1_readdata),   //                    .readdata
		.out_port   (pio_led_external_connection_export)       // external_connection.export
	);

	top_pll_0 pll_0 (
		.refclk   (clk_clk),                  //  refclk.clk
		.rst      (~reset_reset_n),           //   reset.reset
		.outclk_0 (pll_0_outclk0_clk),        // outclk0.clk
		.outclk_1 (pll_0_outclk1_100mhz_clk), // outclk1.clk
		.outclk_2 (pll_0_outclk2_20mhz_clk),  // outclk2.clk
		.locked   ()                          // (terminated)
	);

	top_sdram_vfb sdram_vfb (
		.clk            (pll_0_outclk0_clk),                            //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),              // reset.reset_n
		.az_addr        (mm_interconnect_3_sdram_vfb_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_3_sdram_vfb_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_3_sdram_vfb_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_3_sdram_vfb_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_3_sdram_vfb_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_3_sdram_vfb_s1_write),        //      .write_n
		.za_data        (mm_interconnect_3_sdram_vfb_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_3_sdram_vfb_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_3_sdram_vfb_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_vfb_wire_addr),                          //  wire.export
		.zs_ba          (sdram_vfb_wire_ba),                            //      .export
		.zs_cas_n       (sdram_vfb_wire_cas_n),                         //      .export
		.zs_cke         (sdram_vfb_wire_cke),                           //      .export
		.zs_cs_n        (sdram_vfb_wire_cs_n),                          //      .export
		.zs_dq          (sdram_vfb_wire_dq),                            //      .export
		.zs_dqm         (sdram_vfb_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_vfb_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_vfb_wire_we_n)                           //      .export
	);

	top_sysid_qsys_0 sysid_qsys_0 (
		.clock    (pll_0_outclk0_clk),                                     //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //         reset.reset_n
		.readdata (mm_interconnect_1_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_1_sysid_qsys_0_control_slave_address)   //              .address
	);

	top_timer_0 timer_0 (
		.clk        (pll_0_outclk0_clk),                       //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_1_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver5_irq)                 //   irq.irq
	);

	top_mm_interconnect_0 mm_interconnect_0 (
		.pcie_256_dma_coreclkout_clk                   (pcie_256_dma_coreclkout_clk),                //                 pcie_256_dma_coreclkout.clk
		.csr_regmap_reset2_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),         // csr_regmap_reset2_reset_bridge_in_reset.reset
		.pcie_256_dma_Rxm_BAR2_address                 (pcie_256_dma_rxm_bar2_address),              //                   pcie_256_dma_Rxm_BAR2.address
		.pcie_256_dma_Rxm_BAR2_waitrequest             (pcie_256_dma_rxm_bar2_waitrequest),          //                                        .waitrequest
		.pcie_256_dma_Rxm_BAR2_byteenable              (pcie_256_dma_rxm_bar2_byteenable),           //                                        .byteenable
		.pcie_256_dma_Rxm_BAR2_read                    (pcie_256_dma_rxm_bar2_read),                 //                                        .read
		.pcie_256_dma_Rxm_BAR2_readdata                (pcie_256_dma_rxm_bar2_readdata),             //                                        .readdata
		.pcie_256_dma_Rxm_BAR2_readdatavalid           (pcie_256_dma_rxm_bar2_readdatavalid),        //                                        .readdatavalid
		.pcie_256_dma_Rxm_BAR2_write                   (pcie_256_dma_rxm_bar2_write),                //                                        .write
		.pcie_256_dma_Rxm_BAR2_writedata               (pcie_256_dma_rxm_bar2_writedata),            //                                        .writedata
		.csr_regmap_s2_address                         (mm_interconnect_0_csr_regmap_s2_address),    //                           csr_regmap_s2.address
		.csr_regmap_s2_write                           (mm_interconnect_0_csr_regmap_s2_write),      //                                        .write
		.csr_regmap_s2_readdata                        (mm_interconnect_0_csr_regmap_s2_readdata),   //                                        .readdata
		.csr_regmap_s2_writedata                       (mm_interconnect_0_csr_regmap_s2_writedata),  //                                        .writedata
		.csr_regmap_s2_byteenable                      (mm_interconnect_0_csr_regmap_s2_byteenable), //                                        .byteenable
		.csr_regmap_s2_chipselect                      (mm_interconnect_0_csr_regmap_s2_chipselect), //                                        .chipselect
		.csr_regmap_s2_clken                           (mm_interconnect_0_csr_regmap_s2_clken)       //                                        .clken
	);

	top_mm_interconnect_1 mm_interconnect_1 (
		.pll_0_outclk0_clk                                               (pll_0_outclk0_clk),                                                  //                                             pll_0_outclk0.clk
		.mem_if_ddr3_emif_0_mp_cmd_reset_n_0_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                     // mem_if_ddr3_emif_0_mp_cmd_reset_n_0_reset_bridge_in_reset.reset
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset                  (rst_controller_reset_out_reset),                                     //                  nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address                                (nios2_gen2_0_data_master_address),                                   //                                  nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest                            (nios2_gen2_0_data_master_waitrequest),                               //                                                          .waitrequest
		.nios2_gen2_0_data_master_byteenable                             (nios2_gen2_0_data_master_byteenable),                                //                                                          .byteenable
		.nios2_gen2_0_data_master_read                                   (nios2_gen2_0_data_master_read),                                      //                                                          .read
		.nios2_gen2_0_data_master_readdata                               (nios2_gen2_0_data_master_readdata),                                  //                                                          .readdata
		.nios2_gen2_0_data_master_readdatavalid                          (nios2_gen2_0_data_master_readdatavalid),                             //                                                          .readdatavalid
		.nios2_gen2_0_data_master_write                                  (nios2_gen2_0_data_master_write),                                     //                                                          .write
		.nios2_gen2_0_data_master_writedata                              (nios2_gen2_0_data_master_writedata),                                 //                                                          .writedata
		.nios2_gen2_0_data_master_debugaccess                            (nios2_gen2_0_data_master_debugaccess),                               //                                                          .debugaccess
		.nios2_gen2_0_instruction_master_address                         (nios2_gen2_0_instruction_master_address),                            //                           nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest                     (nios2_gen2_0_instruction_master_waitrequest),                        //                                                          .waitrequest
		.nios2_gen2_0_instruction_master_read                            (nios2_gen2_0_instruction_master_read),                               //                                                          .read
		.nios2_gen2_0_instruction_master_readdata                        (nios2_gen2_0_instruction_master_readdata),                           //                                                          .readdata
		.nios2_gen2_0_instruction_master_readdatavalid                   (nios2_gen2_0_instruction_master_readdatavalid),                      //                                                          .readdatavalid
		.csr_regmap_s1_address                                           (mm_interconnect_1_csr_regmap_s1_address),                            //                                             csr_regmap_s1.address
		.csr_regmap_s1_write                                             (mm_interconnect_1_csr_regmap_s1_write),                              //                                                          .write
		.csr_regmap_s1_readdata                                          (mm_interconnect_1_csr_regmap_s1_readdata),                           //                                                          .readdata
		.csr_regmap_s1_writedata                                         (mm_interconnect_1_csr_regmap_s1_writedata),                          //                                                          .writedata
		.csr_regmap_s1_byteenable                                        (mm_interconnect_1_csr_regmap_s1_byteenable),                         //                                                          .byteenable
		.csr_regmap_s1_chipselect                                        (mm_interconnect_1_csr_regmap_s1_chipselect),                         //                                                          .chipselect
		.csr_regmap_s1_clken                                             (mm_interconnect_1_csr_regmap_s1_clken),                              //                                                          .clken
		.ddr3_status_s1_address                                          (mm_interconnect_1_ddr3_status_s1_address),                           //                                            ddr3_status_s1.address
		.ddr3_status_s1_readdata                                         (mm_interconnect_1_ddr3_status_s1_readdata),                          //                                                          .readdata
		.fifo_0_in_csr_address                                           (mm_interconnect_1_fifo_0_in_csr_address),                            //                                             fifo_0_in_csr.address
		.fifo_0_in_csr_write                                             (mm_interconnect_1_fifo_0_in_csr_write),                              //                                                          .write
		.fifo_0_in_csr_read                                              (mm_interconnect_1_fifo_0_in_csr_read),                               //                                                          .read
		.fifo_0_in_csr_readdata                                          (mm_interconnect_1_fifo_0_in_csr_readdata),                           //                                                          .readdata
		.fifo_0_in_csr_writedata                                         (mm_interconnect_1_fifo_0_in_csr_writedata),                          //                                                          .writedata
		.fifo_0_out_address                                              (mm_interconnect_1_fifo_0_out_address),                               //                                                fifo_0_out.address
		.fifo_0_out_read                                                 (mm_interconnect_1_fifo_0_out_read),                                  //                                                          .read
		.fifo_0_out_readdata                                             (mm_interconnect_1_fifo_0_out_readdata),                              //                                                          .readdata
		.fifo_0_out_waitrequest                                          (mm_interconnect_1_fifo_0_out_waitrequest),                           //                                                          .waitrequest
		.i2c_opencores_camera_avalon_slave_0_address                     (mm_interconnect_1_i2c_opencores_camera_avalon_slave_0_address),      //                       i2c_opencores_camera_avalon_slave_0.address
		.i2c_opencores_camera_avalon_slave_0_write                       (mm_interconnect_1_i2c_opencores_camera_avalon_slave_0_write),        //                                                          .write
		.i2c_opencores_camera_avalon_slave_0_readdata                    (mm_interconnect_1_i2c_opencores_camera_avalon_slave_0_readdata),     //                                                          .readdata
		.i2c_opencores_camera_avalon_slave_0_writedata                   (mm_interconnect_1_i2c_opencores_camera_avalon_slave_0_writedata),    //                                                          .writedata
		.i2c_opencores_camera_avalon_slave_0_waitrequest                 (~mm_interconnect_1_i2c_opencores_camera_avalon_slave_0_waitrequest), //                                                          .waitrequest
		.i2c_opencores_camera_avalon_slave_0_chipselect                  (mm_interconnect_1_i2c_opencores_camera_avalon_slave_0_chipselect),   //                                                          .chipselect
		.i2c_opencores_mipi_avalon_slave_0_address                       (mm_interconnect_1_i2c_opencores_mipi_avalon_slave_0_address),        //                         i2c_opencores_mipi_avalon_slave_0.address
		.i2c_opencores_mipi_avalon_slave_0_write                         (mm_interconnect_1_i2c_opencores_mipi_avalon_slave_0_write),          //                                                          .write
		.i2c_opencores_mipi_avalon_slave_0_readdata                      (mm_interconnect_1_i2c_opencores_mipi_avalon_slave_0_readdata),       //                                                          .readdata
		.i2c_opencores_mipi_avalon_slave_0_writedata                     (mm_interconnect_1_i2c_opencores_mipi_avalon_slave_0_writedata),      //                                                          .writedata
		.i2c_opencores_mipi_avalon_slave_0_waitrequest                   (~mm_interconnect_1_i2c_opencores_mipi_avalon_slave_0_waitrequest),   //                                                          .waitrequest
		.i2c_opencores_mipi_avalon_slave_0_chipselect                    (mm_interconnect_1_i2c_opencores_mipi_avalon_slave_0_chipselect),     //                                                          .chipselect
		.jtag_uart_0_avalon_jtag_slave_address                           (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_address),            //                             jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write                             (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write),              //                                                          .write
		.jtag_uart_0_avalon_jtag_slave_read                              (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read),               //                                                          .read
		.jtag_uart_0_avalon_jtag_slave_readdata                          (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_readdata),           //                                                          .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata                         (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_writedata),          //                                                          .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest                       (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_waitrequest),        //                                                          .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect                        (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_chipselect),         //                                                          .chipselect
		.mem_if_ddr3_emif_0_avl_0_address                                (mm_interconnect_1_mem_if_ddr3_emif_0_avl_0_address),                 //                                  mem_if_ddr3_emif_0_avl_0.address
		.mem_if_ddr3_emif_0_avl_0_write                                  (mm_interconnect_1_mem_if_ddr3_emif_0_avl_0_write),                   //                                                          .write
		.mem_if_ddr3_emif_0_avl_0_read                                   (mm_interconnect_1_mem_if_ddr3_emif_0_avl_0_read),                    //                                                          .read
		.mem_if_ddr3_emif_0_avl_0_readdata                               (mm_interconnect_1_mem_if_ddr3_emif_0_avl_0_readdata),                //                                                          .readdata
		.mem_if_ddr3_emif_0_avl_0_writedata                              (mm_interconnect_1_mem_if_ddr3_emif_0_avl_0_writedata),               //                                                          .writedata
		.mem_if_ddr3_emif_0_avl_0_beginbursttransfer                     (mm_interconnect_1_mem_if_ddr3_emif_0_avl_0_beginbursttransfer),      //                                                          .beginbursttransfer
		.mem_if_ddr3_emif_0_avl_0_burstcount                             (mm_interconnect_1_mem_if_ddr3_emif_0_avl_0_burstcount),              //                                                          .burstcount
		.mem_if_ddr3_emif_0_avl_0_byteenable                             (mm_interconnect_1_mem_if_ddr3_emif_0_avl_0_byteenable),              //                                                          .byteenable
		.mem_if_ddr3_emif_0_avl_0_readdatavalid                          (mm_interconnect_1_mem_if_ddr3_emif_0_avl_0_readdatavalid),           //                                                          .readdatavalid
		.mem_if_ddr3_emif_0_avl_0_waitrequest                            (~mm_interconnect_1_mem_if_ddr3_emif_0_avl_0_waitrequest),            //                                                          .waitrequest
		.mipi_pwdn_n_s1_address                                          (mm_interconnect_1_mipi_pwdn_n_s1_address),                           //                                            mipi_pwdn_n_s1.address
		.mipi_pwdn_n_s1_write                                            (mm_interconnect_1_mipi_pwdn_n_s1_write),                             //                                                          .write
		.mipi_pwdn_n_s1_readdata                                         (mm_interconnect_1_mipi_pwdn_n_s1_readdata),                          //                                                          .readdata
		.mipi_pwdn_n_s1_writedata                                        (mm_interconnect_1_mipi_pwdn_n_s1_writedata),                         //                                                          .writedata
		.mipi_pwdn_n_s1_chipselect                                       (mm_interconnect_1_mipi_pwdn_n_s1_chipselect),                        //                                                          .chipselect
		.mipi_reset_n_s1_address                                         (mm_interconnect_1_mipi_reset_n_s1_address),                          //                                           mipi_reset_n_s1.address
		.mipi_reset_n_s1_write                                           (mm_interconnect_1_mipi_reset_n_s1_write),                            //                                                          .write
		.mipi_reset_n_s1_readdata                                        (mm_interconnect_1_mipi_reset_n_s1_readdata),                         //                                                          .readdata
		.mipi_reset_n_s1_writedata                                       (mm_interconnect_1_mipi_reset_n_s1_writedata),                        //                                                          .writedata
		.mipi_reset_n_s1_chipselect                                      (mm_interconnect_1_mipi_reset_n_s1_chipselect),                       //                                                          .chipselect
		.nios2_gen2_0_debug_mem_slave_address                            (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_address),             //                              nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write                              (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_write),               //                                                          .write
		.nios2_gen2_0_debug_mem_slave_read                               (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_read),                //                                                          .read
		.nios2_gen2_0_debug_mem_slave_readdata                           (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_readdata),            //                                                          .readdata
		.nios2_gen2_0_debug_mem_slave_writedata                          (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_writedata),           //                                                          .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable                         (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_byteenable),          //                                                          .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest                        (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_waitrequest),         //                                                          .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess                        (mm_interconnect_1_nios2_gen2_0_debug_mem_slave_debugaccess),         //                                                          .debugaccess
		.nios_ram_s1_address                                             (mm_interconnect_1_nios_ram_s1_address),                              //                                               nios_ram_s1.address
		.nios_ram_s1_write                                               (mm_interconnect_1_nios_ram_s1_write),                                //                                                          .write
		.nios_ram_s1_readdata                                            (mm_interconnect_1_nios_ram_s1_readdata),                             //                                                          .readdata
		.nios_ram_s1_writedata                                           (mm_interconnect_1_nios_ram_s1_writedata),                            //                                                          .writedata
		.nios_ram_s1_byteenable                                          (mm_interconnect_1_nios_ram_s1_byteenable),                           //                                                          .byteenable
		.nios_ram_s1_chipselect                                          (mm_interconnect_1_nios_ram_s1_chipselect),                           //                                                          .chipselect
		.nios_ram_s1_clken                                               (mm_interconnect_1_nios_ram_s1_clken),                                //                                                          .clken
		.ocm_256k_dma_s1_address                                         (mm_interconnect_1_ocm_256k_dma_s1_address),                          //                                           ocm_256k_dma_s1.address
		.ocm_256k_dma_s1_write                                           (mm_interconnect_1_ocm_256k_dma_s1_write),                            //                                                          .write
		.ocm_256k_dma_s1_readdata                                        (mm_interconnect_1_ocm_256k_dma_s1_readdata),                         //                                                          .readdata
		.ocm_256k_dma_s1_writedata                                       (mm_interconnect_1_ocm_256k_dma_s1_writedata),                        //                                                          .writedata
		.ocm_256k_dma_s1_byteenable                                      (mm_interconnect_1_ocm_256k_dma_s1_byteenable),                       //                                                          .byteenable
		.ocm_256k_dma_s1_chipselect                                      (mm_interconnect_1_ocm_256k_dma_s1_chipselect),                       //                                                          .chipselect
		.ocm_256k_dma_s1_clken                                           (mm_interconnect_1_ocm_256k_dma_s1_clken),                            //                                                          .clken
		.pio_button_s1_address                                           (mm_interconnect_1_pio_button_s1_address),                            //                                             pio_button_s1.address
		.pio_button_s1_write                                             (mm_interconnect_1_pio_button_s1_write),                              //                                                          .write
		.pio_button_s1_readdata                                          (mm_interconnect_1_pio_button_s1_readdata),                           //                                                          .readdata
		.pio_button_s1_writedata                                         (mm_interconnect_1_pio_button_s1_writedata),                          //                                                          .writedata
		.pio_button_s1_chipselect                                        (mm_interconnect_1_pio_button_s1_chipselect),                         //                                                          .chipselect
		.pio_led_s1_address                                              (mm_interconnect_1_pio_led_s1_address),                               //                                                pio_led_s1.address
		.pio_led_s1_write                                                (mm_interconnect_1_pio_led_s1_write),                                 //                                                          .write
		.pio_led_s1_readdata                                             (mm_interconnect_1_pio_led_s1_readdata),                              //                                                          .readdata
		.pio_led_s1_writedata                                            (mm_interconnect_1_pio_led_s1_writedata),                             //                                                          .writedata
		.pio_led_s1_chipselect                                           (mm_interconnect_1_pio_led_s1_chipselect),                            //                                                          .chipselect
		.sysid_qsys_0_control_slave_address                              (mm_interconnect_1_sysid_qsys_0_control_slave_address),               //                                sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata                             (mm_interconnect_1_sysid_qsys_0_control_slave_readdata),              //                                                          .readdata
		.TERASIC_AUTO_FOCUS_0_mm_ctrl_address                            (mm_interconnect_1_terasic_auto_focus_0_mm_ctrl_address),             //                              TERASIC_AUTO_FOCUS_0_mm_ctrl.address
		.TERASIC_AUTO_FOCUS_0_mm_ctrl_write                              (mm_interconnect_1_terasic_auto_focus_0_mm_ctrl_write),               //                                                          .write
		.TERASIC_AUTO_FOCUS_0_mm_ctrl_read                               (mm_interconnect_1_terasic_auto_focus_0_mm_ctrl_read),                //                                                          .read
		.TERASIC_AUTO_FOCUS_0_mm_ctrl_readdata                           (mm_interconnect_1_terasic_auto_focus_0_mm_ctrl_readdata),            //                                                          .readdata
		.TERASIC_AUTO_FOCUS_0_mm_ctrl_writedata                          (mm_interconnect_1_terasic_auto_focus_0_mm_ctrl_writedata),           //                                                          .writedata
		.TERASIC_AUTO_FOCUS_0_mm_ctrl_chipselect                         (mm_interconnect_1_terasic_auto_focus_0_mm_ctrl_chipselect),          //                                                          .chipselect
		.timer_0_s1_address                                              (mm_interconnect_1_timer_0_s1_address),                               //                                                timer_0_s1.address
		.timer_0_s1_write                                                (mm_interconnect_1_timer_0_s1_write),                                 //                                                          .write
		.timer_0_s1_readdata                                             (mm_interconnect_1_timer_0_s1_readdata),                              //                                                          .readdata
		.timer_0_s1_writedata                                            (mm_interconnect_1_timer_0_s1_writedata),                             //                                                          .writedata
		.timer_0_s1_chipselect                                           (mm_interconnect_1_timer_0_s1_chipselect)                             //                                                          .chipselect
	);

	top_mm_interconnect_2 mm_interconnect_2 (
		.pcie_256_dma_coreclkout_clk                     (pcie_256_dma_coreclkout_clk),                             //                   pcie_256_dma_coreclkout.clk
		.ocm_256k_dma_reset2_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                      // ocm_256k_dma_reset2_reset_bridge_in_reset.reset
		.pcie_256_dma_dma_rd_master_address              (pcie_256_dma_dma_rd_master_address),                      //                pcie_256_dma_dma_rd_master.address
		.pcie_256_dma_dma_rd_master_waitrequest          (pcie_256_dma_dma_rd_master_waitrequest),                  //                                          .waitrequest
		.pcie_256_dma_dma_rd_master_burstcount           (pcie_256_dma_dma_rd_master_burstcount),                   //                                          .burstcount
		.pcie_256_dma_dma_rd_master_byteenable           (pcie_256_dma_dma_rd_master_byteenable),                   //                                          .byteenable
		.pcie_256_dma_dma_rd_master_write                (pcie_256_dma_dma_rd_master_write),                        //                                          .write
		.pcie_256_dma_dma_rd_master_writedata            (pcie_256_dma_dma_rd_master_writedata),                    //                                          .writedata
		.pcie_256_dma_dma_wr_master_address              (pcie_256_dma_dma_wr_master_address),                      //                pcie_256_dma_dma_wr_master.address
		.pcie_256_dma_dma_wr_master_waitrequest          (pcie_256_dma_dma_wr_master_waitrequest),                  //                                          .waitrequest
		.pcie_256_dma_dma_wr_master_burstcount           (pcie_256_dma_dma_wr_master_burstcount),                   //                                          .burstcount
		.pcie_256_dma_dma_wr_master_read                 (pcie_256_dma_dma_wr_master_read),                         //                                          .read
		.pcie_256_dma_dma_wr_master_readdata             (pcie_256_dma_dma_wr_master_readdata),                     //                                          .readdata
		.pcie_256_dma_dma_wr_master_readdatavalid        (pcie_256_dma_dma_wr_master_readdatavalid),                //                                          .readdatavalid
		.ocm_256k_dma_s2_address                         (mm_interconnect_2_ocm_256k_dma_s2_address),               //                           ocm_256k_dma_s2.address
		.ocm_256k_dma_s2_write                           (mm_interconnect_2_ocm_256k_dma_s2_write),                 //                                          .write
		.ocm_256k_dma_s2_readdata                        (mm_interconnect_2_ocm_256k_dma_s2_readdata),              //                                          .readdata
		.ocm_256k_dma_s2_writedata                       (mm_interconnect_2_ocm_256k_dma_s2_writedata),             //                                          .writedata
		.ocm_256k_dma_s2_byteenable                      (mm_interconnect_2_ocm_256k_dma_s2_byteenable),            //                                          .byteenable
		.ocm_256k_dma_s2_chipselect                      (mm_interconnect_2_ocm_256k_dma_s2_chipselect),            //                                          .chipselect
		.ocm_256k_dma_s2_clken                           (mm_interconnect_2_ocm_256k_dma_s2_clken),                 //                                          .clken
		.pcie_256_dma_rd_dts_slave_address               (mm_interconnect_2_pcie_256_dma_rd_dts_slave_address),     //                 pcie_256_dma_rd_dts_slave.address
		.pcie_256_dma_rd_dts_slave_write                 (mm_interconnect_2_pcie_256_dma_rd_dts_slave_write),       //                                          .write
		.pcie_256_dma_rd_dts_slave_writedata             (mm_interconnect_2_pcie_256_dma_rd_dts_slave_writedata),   //                                          .writedata
		.pcie_256_dma_rd_dts_slave_burstcount            (mm_interconnect_2_pcie_256_dma_rd_dts_slave_burstcount),  //                                          .burstcount
		.pcie_256_dma_rd_dts_slave_waitrequest           (mm_interconnect_2_pcie_256_dma_rd_dts_slave_waitrequest), //                                          .waitrequest
		.pcie_256_dma_rd_dts_slave_chipselect            (mm_interconnect_2_pcie_256_dma_rd_dts_slave_chipselect),  //                                          .chipselect
		.pcie_256_dma_wr_dts_slave_address               (mm_interconnect_2_pcie_256_dma_wr_dts_slave_address),     //                 pcie_256_dma_wr_dts_slave.address
		.pcie_256_dma_wr_dts_slave_write                 (mm_interconnect_2_pcie_256_dma_wr_dts_slave_write),       //                                          .write
		.pcie_256_dma_wr_dts_slave_writedata             (mm_interconnect_2_pcie_256_dma_wr_dts_slave_writedata),   //                                          .writedata
		.pcie_256_dma_wr_dts_slave_burstcount            (mm_interconnect_2_pcie_256_dma_wr_dts_slave_burstcount),  //                                          .burstcount
		.pcie_256_dma_wr_dts_slave_waitrequest           (mm_interconnect_2_pcie_256_dma_wr_dts_slave_waitrequest), //                                          .waitrequest
		.pcie_256_dma_wr_dts_slave_chipselect            (mm_interconnect_2_pcie_256_dma_wr_dts_slave_chipselect)   //                                          .chipselect
	);

	top_mm_interconnect_3 mm_interconnect_3 (
		.pll_0_outclk0_clk                                       (pll_0_outclk0_clk),                            //                                     pll_0_outclk0.clk
		.alt_vip_cl_vfb_0_main_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),               // alt_vip_cl_vfb_0_main_reset_reset_bridge_in_reset.reset
		.alt_vip_cl_vfb_0_mem_master_rd_address                  (alt_vip_cl_vfb_0_mem_master_rd_address),       //                    alt_vip_cl_vfb_0_mem_master_rd.address
		.alt_vip_cl_vfb_0_mem_master_rd_waitrequest              (alt_vip_cl_vfb_0_mem_master_rd_waitrequest),   //                                                  .waitrequest
		.alt_vip_cl_vfb_0_mem_master_rd_burstcount               (alt_vip_cl_vfb_0_mem_master_rd_burstcount),    //                                                  .burstcount
		.alt_vip_cl_vfb_0_mem_master_rd_read                     (alt_vip_cl_vfb_0_mem_master_rd_read),          //                                                  .read
		.alt_vip_cl_vfb_0_mem_master_rd_readdata                 (alt_vip_cl_vfb_0_mem_master_rd_readdata),      //                                                  .readdata
		.alt_vip_cl_vfb_0_mem_master_rd_readdatavalid            (alt_vip_cl_vfb_0_mem_master_rd_readdatavalid), //                                                  .readdatavalid
		.alt_vip_cl_vfb_0_mem_master_wr_address                  (alt_vip_cl_vfb_0_mem_master_wr_address),       //                    alt_vip_cl_vfb_0_mem_master_wr.address
		.alt_vip_cl_vfb_0_mem_master_wr_waitrequest              (alt_vip_cl_vfb_0_mem_master_wr_waitrequest),   //                                                  .waitrequest
		.alt_vip_cl_vfb_0_mem_master_wr_burstcount               (alt_vip_cl_vfb_0_mem_master_wr_burstcount),    //                                                  .burstcount
		.alt_vip_cl_vfb_0_mem_master_wr_byteenable               (alt_vip_cl_vfb_0_mem_master_wr_byteenable),    //                                                  .byteenable
		.alt_vip_cl_vfb_0_mem_master_wr_write                    (alt_vip_cl_vfb_0_mem_master_wr_write),         //                                                  .write
		.alt_vip_cl_vfb_0_mem_master_wr_writedata                (alt_vip_cl_vfb_0_mem_master_wr_writedata),     //                                                  .writedata
		.sdram_vfb_s1_address                                    (mm_interconnect_3_sdram_vfb_s1_address),       //                                      sdram_vfb_s1.address
		.sdram_vfb_s1_write                                      (mm_interconnect_3_sdram_vfb_s1_write),         //                                                  .write
		.sdram_vfb_s1_read                                       (mm_interconnect_3_sdram_vfb_s1_read),          //                                                  .read
		.sdram_vfb_s1_readdata                                   (mm_interconnect_3_sdram_vfb_s1_readdata),      //                                                  .readdata
		.sdram_vfb_s1_writedata                                  (mm_interconnect_3_sdram_vfb_s1_writedata),     //                                                  .writedata
		.sdram_vfb_s1_byteenable                                 (mm_interconnect_3_sdram_vfb_s1_byteenable),    //                                                  .byteenable
		.sdram_vfb_s1_readdatavalid                              (mm_interconnect_3_sdram_vfb_s1_readdatavalid), //                                                  .readdatavalid
		.sdram_vfb_s1_waitrequest                                (mm_interconnect_3_sdram_vfb_s1_waitrequest),   //                                                  .waitrequest
		.sdram_vfb_s1_chipselect                                 (mm_interconnect_3_sdram_vfb_s1_chipselect)     //                                                  .chipselect
	);

	top_mm_interconnect_4 mm_interconnect_4 (
		.pcie_256_dma_coreclkout_clk                                             (pcie_256_dma_coreclkout_clk),                      //                                           pcie_256_dma_coreclkout.clk
		.pcie_256_dma_rd_dcm_master_translator_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),               // pcie_256_dma_rd_dcm_master_translator_reset_reset_bridge_in_reset.reset
		.pcie_256_dma_rd_dcm_master_address                                      (pcie_256_dma_rd_dcm_master_address),               //                                        pcie_256_dma_rd_dcm_master.address
		.pcie_256_dma_rd_dcm_master_waitrequest                                  (pcie_256_dma_rd_dcm_master_waitrequest),           //                                                                  .waitrequest
		.pcie_256_dma_rd_dcm_master_byteenable                                   (pcie_256_dma_rd_dcm_master_byteenable),            //                                                                  .byteenable
		.pcie_256_dma_rd_dcm_master_read                                         (pcie_256_dma_rd_dcm_master_read),                  //                                                                  .read
		.pcie_256_dma_rd_dcm_master_readdata                                     (pcie_256_dma_rd_dcm_master_readdata),              //                                                                  .readdata
		.pcie_256_dma_rd_dcm_master_readdatavalid                                (pcie_256_dma_rd_dcm_master_readdatavalid),         //                                                                  .readdatavalid
		.pcie_256_dma_rd_dcm_master_write                                        (pcie_256_dma_rd_dcm_master_write),                 //                                                                  .write
		.pcie_256_dma_rd_dcm_master_writedata                                    (pcie_256_dma_rd_dcm_master_writedata),             //                                                                  .writedata
		.pcie_256_dma_wr_dcm_master_address                                      (pcie_256_dma_wr_dcm_master_address),               //                                        pcie_256_dma_wr_dcm_master.address
		.pcie_256_dma_wr_dcm_master_waitrequest                                  (pcie_256_dma_wr_dcm_master_waitrequest),           //                                                                  .waitrequest
		.pcie_256_dma_wr_dcm_master_byteenable                                   (pcie_256_dma_wr_dcm_master_byteenable),            //                                                                  .byteenable
		.pcie_256_dma_wr_dcm_master_read                                         (pcie_256_dma_wr_dcm_master_read),                  //                                                                  .read
		.pcie_256_dma_wr_dcm_master_readdata                                     (pcie_256_dma_wr_dcm_master_readdata),              //                                                                  .readdata
		.pcie_256_dma_wr_dcm_master_readdatavalid                                (pcie_256_dma_wr_dcm_master_readdatavalid),         //                                                                  .readdatavalid
		.pcie_256_dma_wr_dcm_master_write                                        (pcie_256_dma_wr_dcm_master_write),                 //                                                                  .write
		.pcie_256_dma_wr_dcm_master_writedata                                    (pcie_256_dma_wr_dcm_master_writedata),             //                                                                  .writedata
		.pcie_256_dma_Txs_address                                                (mm_interconnect_4_pcie_256_dma_txs_address),       //                                                  pcie_256_dma_Txs.address
		.pcie_256_dma_Txs_write                                                  (mm_interconnect_4_pcie_256_dma_txs_write),         //                                                                  .write
		.pcie_256_dma_Txs_read                                                   (mm_interconnect_4_pcie_256_dma_txs_read),          //                                                                  .read
		.pcie_256_dma_Txs_readdata                                               (mm_interconnect_4_pcie_256_dma_txs_readdata),      //                                                                  .readdata
		.pcie_256_dma_Txs_writedata                                              (mm_interconnect_4_pcie_256_dma_txs_writedata),     //                                                                  .writedata
		.pcie_256_dma_Txs_byteenable                                             (mm_interconnect_4_pcie_256_dma_txs_byteenable),    //                                                                  .byteenable
		.pcie_256_dma_Txs_readdatavalid                                          (mm_interconnect_4_pcie_256_dma_txs_readdatavalid), //                                                                  .readdatavalid
		.pcie_256_dma_Txs_waitrequest                                            (mm_interconnect_4_pcie_256_dma_txs_waitrequest),   //                                                                  .waitrequest
		.pcie_256_dma_Txs_chipselect                                             (mm_interconnect_4_pcie_256_dma_txs_chipselect)     //                                                                  .chipselect
	);

	top_mm_interconnect_5 mm_interconnect_5 (
		.clk_0_clk_clk                                                        (clk_clk),                                                         //                                                      clk_0_clk.clk
		.pcie_256_dma_coreclkout_clk                                          (pcie_256_dma_coreclkout_clk),                                     //                                        pcie_256_dma_coreclkout.clk
		.alt_xcvr_reconfig_0_mgmt_rst_reset_reset_bridge_in_reset_reset       (rst_controller_001_reset_out_reset),                              //       alt_xcvr_reconfig_0_mgmt_rst_reset_reset_bridge_in_reset.reset
		.pcie_reconfig_driver_0_reconfig_xcvr_rst_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                              // pcie_reconfig_driver_0_reconfig_xcvr_rst_reset_bridge_in_reset.reset
		.pcie_reconfig_driver_0_reconfig_mgmt_address                         (pcie_reconfig_driver_0_reconfig_mgmt_address),                    //                           pcie_reconfig_driver_0_reconfig_mgmt.address
		.pcie_reconfig_driver_0_reconfig_mgmt_waitrequest                     (pcie_reconfig_driver_0_reconfig_mgmt_waitrequest),                //                                                               .waitrequest
		.pcie_reconfig_driver_0_reconfig_mgmt_read                            (pcie_reconfig_driver_0_reconfig_mgmt_read),                       //                                                               .read
		.pcie_reconfig_driver_0_reconfig_mgmt_readdata                        (pcie_reconfig_driver_0_reconfig_mgmt_readdata),                   //                                                               .readdata
		.pcie_reconfig_driver_0_reconfig_mgmt_write                           (pcie_reconfig_driver_0_reconfig_mgmt_write),                      //                                                               .write
		.pcie_reconfig_driver_0_reconfig_mgmt_writedata                       (pcie_reconfig_driver_0_reconfig_mgmt_writedata),                  //                                                               .writedata
		.alt_xcvr_reconfig_0_reconfig_mgmt_address                            (mm_interconnect_5_alt_xcvr_reconfig_0_reconfig_mgmt_address),     //                              alt_xcvr_reconfig_0_reconfig_mgmt.address
		.alt_xcvr_reconfig_0_reconfig_mgmt_write                              (mm_interconnect_5_alt_xcvr_reconfig_0_reconfig_mgmt_write),       //                                                               .write
		.alt_xcvr_reconfig_0_reconfig_mgmt_read                               (mm_interconnect_5_alt_xcvr_reconfig_0_reconfig_mgmt_read),        //                                                               .read
		.alt_xcvr_reconfig_0_reconfig_mgmt_readdata                           (mm_interconnect_5_alt_xcvr_reconfig_0_reconfig_mgmt_readdata),    //                                                               .readdata
		.alt_xcvr_reconfig_0_reconfig_mgmt_writedata                          (mm_interconnect_5_alt_xcvr_reconfig_0_reconfig_mgmt_writedata),   //                                                               .writedata
		.alt_xcvr_reconfig_0_reconfig_mgmt_waitrequest                        (mm_interconnect_5_alt_xcvr_reconfig_0_reconfig_mgmt_waitrequest)  //                                                               .waitrequest
	);

	top_irq_mapper irq_mapper (
		.clk           (pll_0_outclk0_clk),              //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),       // receiver5.irq
		.sender_irq    (nios2_gen2_0_irq_irq)            //    sender.irq
	);

	top_avalon_st_adapter #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (24),
		.inChannelWidth  (0),
		.inErrorWidth    (0),
		.inUseEmptyPort  (0),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (24),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (0),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (1)
	) avalon_st_adapter (
		.in_clk_0_clk        (pll_0_outclk0_clk),                                      // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),                         // in_rst_0.reset
		.in_0_data           (terasic_camera_0_avalon_streaming_source_data),          //     in_0.data
		.in_0_valid          (terasic_camera_0_avalon_streaming_source_valid),         //         .valid
		.in_0_ready          (terasic_camera_0_avalon_streaming_source_ready),         //         .ready
		.in_0_startofpacket  (terasic_camera_0_avalon_streaming_source_startofpacket), //         .startofpacket
		.in_0_endofpacket    (terasic_camera_0_avalon_streaming_source_endofpacket),   //         .endofpacket
		.out_0_data          (avalon_st_adapter_out_0_data),                           //    out_0.data
		.out_0_valid         (avalon_st_adapter_out_0_valid),                          //         .valid
		.out_0_ready         (avalon_st_adapter_out_0_ready),                          //         .ready
		.out_0_startofpacket (avalon_st_adapter_out_0_startofpacket),                  //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_out_0_endofpacket)                     //         .endofpacket
	);

	top_avalon_st_adapter_001 #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (32),
		.inChannelWidth  (0),
		.inErrorWidth    (0),
		.inUseEmptyPort  (0),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (1),
		.outDataWidth    (32),
		.outChannelWidth (8),
		.outErrorWidth   (8),
		.outUseEmptyPort (1),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (1)
	) avalon_st_adapter_001 (
		.in_clk_0_clk        (pll_0_outclk0_clk),                         // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),            // in_rst_0.reset
		.in_0_data           (terasic_auto_focus_0_dout_data),            //     in_0.data
		.in_0_valid          (terasic_auto_focus_0_dout_valid),           //         .valid
		.in_0_ready          (terasic_auto_focus_0_dout_ready),           //         .ready
		.in_0_startofpacket  (terasic_auto_focus_0_dout_startofpacket),   //         .startofpacket
		.in_0_endofpacket    (terasic_auto_focus_0_dout_endofpacket),     //         .endofpacket
		.out_0_data          (avalon_st_adapter_001_out_0_data),          //    out_0.data
		.out_0_valid         (avalon_st_adapter_001_out_0_valid),         //         .valid
		.out_0_ready         (avalon_st_adapter_001_out_0_ready),         //         .ready
		.out_0_startofpacket (avalon_st_adapter_001_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_001_out_0_endofpacket),   //         .endofpacket
		.out_0_empty         (avalon_st_adapter_001_out_0_empty),         //         .empty
		.out_0_error         (avalon_st_adapter_001_out_0_error),         //         .error
		.out_0_channel       (avalon_st_adapter_001_out_0_channel)        //         .channel
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (pll_0_outclk0_clk),                  //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~pcie_256_dma_nreset_status_reset),      // reset_in0.reset
		.clk            (pcie_256_dma_coreclkout_clk),            //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_002_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
