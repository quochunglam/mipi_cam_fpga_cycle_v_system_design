// c5_niosii_spi_slvsec.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module c5_niosii_spi_slvsec (
		output wire       b_laser_en_b_laser_en_o,   //   b_laser_en.b_laser_en_o
		input  wire       clk_clk,                   //          clk.clk
		output wire       dlp_en_o_dlp_en_o,         //     dlp_en_o.dlp_en_o
		output wire       inck_en_inck_en_o,         //      inck_en.inck_en_o
		input  wire       key_export,                //          key.export
		output wire [7:0] led_export,                //          led.export
		output wire       r_laser_en_o_r_laser_en_o, // r_laser_en_o.r_laser_en_o
		output wire       reg_1v2_en_reg_1v2_en_o,   //   reg_1v2_en.reg_1v2_en_o
		output wire       reg_1v8_en_reg_1v8_en_o,   //   reg_1v8_en.reg_1v8_en_o
		output wire       reg_3v3_en_reg_3v3_en_o,   //   reg_3v3_en.reg_3v3_en_o
		input  wire       reset_reset_n,             //        reset.reset_n
		input  wire       spi_MISO,                  //          spi.MISO
		output wire       spi_MOSI,                  //             .MOSI
		output wire       spi_SCLK,                  //             .SCLK
		output wire       spi_SS_n,                  //             .SS_n
		input  wire [3:0] sw_export,                 //           sw.export
		output wire       xclr_xclr_o,               //         xclr.xclr_o
		output wire       xtrig_o_xtrig_o            //      xtrig_o.xtrig_o
	);

	wire         pll_0_outclk0_clk;                                              // pll_0:outclk_0 -> [imx421_poweron_0:ctrl_clk_i, laser_dlp_xtrig_controller_0:slave_clk, mm_interconnect_0:pll_0_outclk0_clk, mm_interconnect_1:pll_0_outclk0_clk, niosii_cpu:clk_clk, rst_controller:clk, spi:clk]
	wire         pll_0_outclk1_clk;                                              // pll_0:outclk_1 -> laser_dlp_xtrig_controller_0:ctrl_clk_i
	wire         niosii_cpu_spi_mm_bridge_waitrequest;                           // mm_interconnect_0:niosii_cpu_spi_mm_bridge_waitrequest -> niosii_cpu:spi_mm_bridge_waitrequest
	wire  [31:0] niosii_cpu_spi_mm_bridge_readdata;                              // mm_interconnect_0:niosii_cpu_spi_mm_bridge_readdata -> niosii_cpu:spi_mm_bridge_readdata
	wire         niosii_cpu_spi_mm_bridge_debugaccess;                           // niosii_cpu:spi_mm_bridge_debugaccess -> mm_interconnect_0:niosii_cpu_spi_mm_bridge_debugaccess
	wire   [9:0] niosii_cpu_spi_mm_bridge_address;                               // niosii_cpu:spi_mm_bridge_address -> mm_interconnect_0:niosii_cpu_spi_mm_bridge_address
	wire         niosii_cpu_spi_mm_bridge_read;                                  // niosii_cpu:spi_mm_bridge_read -> mm_interconnect_0:niosii_cpu_spi_mm_bridge_read
	wire   [3:0] niosii_cpu_spi_mm_bridge_byteenable;                            // niosii_cpu:spi_mm_bridge_byteenable -> mm_interconnect_0:niosii_cpu_spi_mm_bridge_byteenable
	wire         niosii_cpu_spi_mm_bridge_readdatavalid;                         // mm_interconnect_0:niosii_cpu_spi_mm_bridge_readdatavalid -> niosii_cpu:spi_mm_bridge_readdatavalid
	wire  [31:0] niosii_cpu_spi_mm_bridge_writedata;                             // niosii_cpu:spi_mm_bridge_writedata -> mm_interconnect_0:niosii_cpu_spi_mm_bridge_writedata
	wire         niosii_cpu_spi_mm_bridge_write;                                 // niosii_cpu:spi_mm_bridge_write -> mm_interconnect_0:niosii_cpu_spi_mm_bridge_write
	wire   [0:0] niosii_cpu_spi_mm_bridge_burstcount;                            // niosii_cpu:spi_mm_bridge_burstcount -> mm_interconnect_0:niosii_cpu_spi_mm_bridge_burstcount
	wire         mm_interconnect_0_spi_spi_control_port_chipselect;              // mm_interconnect_0:spi_spi_control_port_chipselect -> spi:spi_select
	wire  [15:0] mm_interconnect_0_spi_spi_control_port_readdata;                // spi:data_to_cpu -> mm_interconnect_0:spi_spi_control_port_readdata
	wire   [2:0] mm_interconnect_0_spi_spi_control_port_address;                 // mm_interconnect_0:spi_spi_control_port_address -> spi:mem_addr
	wire         mm_interconnect_0_spi_spi_control_port_read;                    // mm_interconnect_0:spi_spi_control_port_read -> spi:read_n
	wire         mm_interconnect_0_spi_spi_control_port_write;                   // mm_interconnect_0:spi_spi_control_port_write -> spi:write_n
	wire  [15:0] mm_interconnect_0_spi_spi_control_port_writedata;               // mm_interconnect_0:spi_spi_control_port_writedata -> spi:data_from_cpu
	wire         niosii_cpu_xtrig_mm_bridge_waitrequest;                         // mm_interconnect_1:niosii_cpu_xtrig_mm_bridge_waitrequest -> niosii_cpu:xtrig_mm_bridge_waitrequest
	wire  [31:0] niosii_cpu_xtrig_mm_bridge_readdata;                            // mm_interconnect_1:niosii_cpu_xtrig_mm_bridge_readdata -> niosii_cpu:xtrig_mm_bridge_readdata
	wire         niosii_cpu_xtrig_mm_bridge_debugaccess;                         // niosii_cpu:xtrig_mm_bridge_debugaccess -> mm_interconnect_1:niosii_cpu_xtrig_mm_bridge_debugaccess
	wire   [9:0] niosii_cpu_xtrig_mm_bridge_address;                             // niosii_cpu:xtrig_mm_bridge_address -> mm_interconnect_1:niosii_cpu_xtrig_mm_bridge_address
	wire         niosii_cpu_xtrig_mm_bridge_read;                                // niosii_cpu:xtrig_mm_bridge_read -> mm_interconnect_1:niosii_cpu_xtrig_mm_bridge_read
	wire   [3:0] niosii_cpu_xtrig_mm_bridge_byteenable;                          // niosii_cpu:xtrig_mm_bridge_byteenable -> mm_interconnect_1:niosii_cpu_xtrig_mm_bridge_byteenable
	wire         niosii_cpu_xtrig_mm_bridge_readdatavalid;                       // mm_interconnect_1:niosii_cpu_xtrig_mm_bridge_readdatavalid -> niosii_cpu:xtrig_mm_bridge_readdatavalid
	wire  [31:0] niosii_cpu_xtrig_mm_bridge_writedata;                           // niosii_cpu:xtrig_mm_bridge_writedata -> mm_interconnect_1:niosii_cpu_xtrig_mm_bridge_writedata
	wire         niosii_cpu_xtrig_mm_bridge_write;                               // niosii_cpu:xtrig_mm_bridge_write -> mm_interconnect_1:niosii_cpu_xtrig_mm_bridge_write
	wire   [0:0] niosii_cpu_xtrig_mm_bridge_burstcount;                          // niosii_cpu:xtrig_mm_bridge_burstcount -> mm_interconnect_1:niosii_cpu_xtrig_mm_bridge_burstcount
	wire  [31:0] mm_interconnect_1_laser_dlp_xtrig_controller_0_avms_readdata;   // laser_dlp_xtrig_controller_0:slave_readdata -> mm_interconnect_1:laser_dlp_xtrig_controller_0_avms_readdata
	wire   [1:0] mm_interconnect_1_laser_dlp_xtrig_controller_0_avms_address;    // mm_interconnect_1:laser_dlp_xtrig_controller_0_avms_address -> laser_dlp_xtrig_controller_0:slave_addr
	wire         mm_interconnect_1_laser_dlp_xtrig_controller_0_avms_read;       // mm_interconnect_1:laser_dlp_xtrig_controller_0_avms_read -> laser_dlp_xtrig_controller_0:slave_read
	wire   [3:0] mm_interconnect_1_laser_dlp_xtrig_controller_0_avms_byteenable; // mm_interconnect_1:laser_dlp_xtrig_controller_0_avms_byteenable -> laser_dlp_xtrig_controller_0:slave_byteenable
	wire         mm_interconnect_1_laser_dlp_xtrig_controller_0_avms_write;      // mm_interconnect_1:laser_dlp_xtrig_controller_0_avms_write -> laser_dlp_xtrig_controller_0:slave_write
	wire  [31:0] mm_interconnect_1_laser_dlp_xtrig_controller_0_avms_writedata;  // mm_interconnect_1:laser_dlp_xtrig_controller_0_avms_writedata -> laser_dlp_xtrig_controller_0:slave_wriredata
	wire         rst_controller_reset_out_reset;                                 // rst_controller:reset_out -> [imx421_poweron_0:ctrl_rst_n_i, mm_interconnect_0:niosii_cpu_reset_reset_bridge_in_reset_reset, mm_interconnect_0:spi_reset_reset_bridge_in_reset_reset, mm_interconnect_1:niosii_cpu_reset_reset_bridge_in_reset_reset, mm_interconnect_1:niosii_cpu_xtrig_mm_bridge_translator_reset_reset_bridge_in_reset_reset, spi:reset_n]

	camera_poweron_sequence_sm #(
		.TIMEOUT_THRESHOLD (34'b0000000000000011110100001001000000)
	) imx421_poweron_0 (
		.ctrl_clk_i   (pll_0_outclk0_clk),               //     clk_in.clk
		.ctrl_rst_n_i (~rst_controller_reset_out_reset), //      rst_n.reset_n
		.reg_1v2_en_o (reg_1v2_en_reg_1v2_en_o),         // reg_1v2_en.reg_1v2_en_o
		.reg_1v8_en_o (reg_1v8_en_reg_1v8_en_o),         // reg_1v8_en.reg_1v8_en_o
		.reg_3v3_en_o (reg_3v3_en_reg_3v3_en_o),         // reg_3v3_en.reg_3v3_en_o
		.inck_en_o    (inck_en_inck_en_o),               //    inck_en.inck_en_o
		.xclr_o       (xclr_xclr_o)                      //       xclr.xclr_o
	);

	laser_dlp_xtrig_controller_avms #(
		.DLP_PULSE_WIDTH (34'b0000000000000000000000000011001000),
		.DATA_WIDTH      (32)
	) laser_dlp_xtrig_controller_0 (
		.slave_addr       (mm_interconnect_1_laser_dlp_xtrig_controller_0_avms_address),    //         avms.address
		.slave_wriredata  (mm_interconnect_1_laser_dlp_xtrig_controller_0_avms_writedata),  //             .writedata
		.slave_byteenable (mm_interconnect_1_laser_dlp_xtrig_controller_0_avms_byteenable), //             .byteenable
		.slave_read       (mm_interconnect_1_laser_dlp_xtrig_controller_0_avms_read),       //             .read
		.slave_readdata   (mm_interconnect_1_laser_dlp_xtrig_controller_0_avms_readdata),   //             .readdata
		.slave_write      (mm_interconnect_1_laser_dlp_xtrig_controller_0_avms_write),      //             .write
		.b_laser_en_o     (b_laser_en_b_laser_en_o),                                        //   b_laser_en.b_laser_en_o
		.r_laser_en_o     (r_laser_en_o_r_laser_en_o),                                      // r_laser_en_o.r_laser_en_o
		.dlp_en_o         (dlp_en_o_dlp_en_o),                                              //     dlp_en_o.dlp_en_o
		.xtrig_o          (xtrig_o_xtrig_o),                                                //      xtrig_o.xtrig_o
		.ctrl_clk_i       (pll_0_outclk1_clk),                                              //          clk.clk
		.ctrl_rst_n_i     (reset_reset_n),                                                  //        rst_n.reset_n
		.slave_clk        (pll_0_outclk0_clk),                                              //     avms_clk.clk
		.slave_reset_n    (reset_reset_n)                                                   //   avms_rst_n.reset_n
	);

	c5_niosii_spi_slvsec_niosii_cpu niosii_cpu (
		.clk_clk                       (pll_0_outclk0_clk),                        //             clk.clk
		.key_export                    (key_export),                               //             key.export
		.led_export                    (led_export),                               //             led.export
		.reset_reset_n                 (reset_reset_n),                            //           reset.reset_n
		.spi_mm_bridge_waitrequest     (niosii_cpu_spi_mm_bridge_waitrequest),     //   spi_mm_bridge.waitrequest
		.spi_mm_bridge_readdata        (niosii_cpu_spi_mm_bridge_readdata),        //                .readdata
		.spi_mm_bridge_readdatavalid   (niosii_cpu_spi_mm_bridge_readdatavalid),   //                .readdatavalid
		.spi_mm_bridge_burstcount      (niosii_cpu_spi_mm_bridge_burstcount),      //                .burstcount
		.spi_mm_bridge_writedata       (niosii_cpu_spi_mm_bridge_writedata),       //                .writedata
		.spi_mm_bridge_address         (niosii_cpu_spi_mm_bridge_address),         //                .address
		.spi_mm_bridge_write           (niosii_cpu_spi_mm_bridge_write),           //                .write
		.spi_mm_bridge_read            (niosii_cpu_spi_mm_bridge_read),            //                .read
		.spi_mm_bridge_byteenable      (niosii_cpu_spi_mm_bridge_byteenable),      //                .byteenable
		.spi_mm_bridge_debugaccess     (niosii_cpu_spi_mm_bridge_debugaccess),     //                .debugaccess
		.sw_export                     (sw_export),                                //              sw.export
		.xtrig_mm_bridge_waitrequest   (niosii_cpu_xtrig_mm_bridge_waitrequest),   // xtrig_mm_bridge.waitrequest
		.xtrig_mm_bridge_readdata      (niosii_cpu_xtrig_mm_bridge_readdata),      //                .readdata
		.xtrig_mm_bridge_readdatavalid (niosii_cpu_xtrig_mm_bridge_readdatavalid), //                .readdatavalid
		.xtrig_mm_bridge_burstcount    (niosii_cpu_xtrig_mm_bridge_burstcount),    //                .burstcount
		.xtrig_mm_bridge_writedata     (niosii_cpu_xtrig_mm_bridge_writedata),     //                .writedata
		.xtrig_mm_bridge_address       (niosii_cpu_xtrig_mm_bridge_address),       //                .address
		.xtrig_mm_bridge_write         (niosii_cpu_xtrig_mm_bridge_write),         //                .write
		.xtrig_mm_bridge_read          (niosii_cpu_xtrig_mm_bridge_read),          //                .read
		.xtrig_mm_bridge_byteenable    (niosii_cpu_xtrig_mm_bridge_byteenable),    //                .byteenable
		.xtrig_mm_bridge_debugaccess   (niosii_cpu_xtrig_mm_bridge_debugaccess)    //                .debugaccess
	);

	c5_niosii_spi_slvsec_pll_0 pll_0 (
		.refclk   (clk_clk),           //  refclk.clk
		.rst      (~reset_reset_n),    //   reset.reset
		.outclk_0 (pll_0_outclk0_clk), // outclk0.clk
		.outclk_1 (pll_0_outclk1_clk), // outclk1.clk
		.locked   ()                   // (terminated)
	);

	c5_niosii_spi_slvsec_spi spi (
		.clk           (pll_0_outclk0_clk),                                 //              clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                   //            reset.reset_n
		.data_from_cpu (mm_interconnect_0_spi_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_0_spi_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_0_spi_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_0_spi_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_0_spi_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_0_spi_spi_control_port_write),     //                 .write_n
		.irq           (),                                                  //              irq.irq
		.MISO          (spi_MISO),                                          //         external.export
		.MOSI          (spi_MOSI),                                          //                 .export
		.SCLK          (spi_SCLK),                                          //                 .export
		.SS_n          (spi_SS_n)                                           //                 .export
	);

	c5_niosii_spi_slvsec_mm_interconnect_0 mm_interconnect_0 (
		.pll_0_outclk0_clk                            (pll_0_outclk0_clk),                                 //                          pll_0_outclk0.clk
		.niosii_cpu_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                    // niosii_cpu_reset_reset_bridge_in_reset.reset
		.spi_reset_reset_bridge_in_reset_reset        (rst_controller_reset_out_reset),                    //        spi_reset_reset_bridge_in_reset.reset
		.niosii_cpu_spi_mm_bridge_address             (niosii_cpu_spi_mm_bridge_address),                  //               niosii_cpu_spi_mm_bridge.address
		.niosii_cpu_spi_mm_bridge_waitrequest         (niosii_cpu_spi_mm_bridge_waitrequest),              //                                       .waitrequest
		.niosii_cpu_spi_mm_bridge_burstcount          (niosii_cpu_spi_mm_bridge_burstcount),               //                                       .burstcount
		.niosii_cpu_spi_mm_bridge_byteenable          (niosii_cpu_spi_mm_bridge_byteenable),               //                                       .byteenable
		.niosii_cpu_spi_mm_bridge_read                (niosii_cpu_spi_mm_bridge_read),                     //                                       .read
		.niosii_cpu_spi_mm_bridge_readdata            (niosii_cpu_spi_mm_bridge_readdata),                 //                                       .readdata
		.niosii_cpu_spi_mm_bridge_readdatavalid       (niosii_cpu_spi_mm_bridge_readdatavalid),            //                                       .readdatavalid
		.niosii_cpu_spi_mm_bridge_write               (niosii_cpu_spi_mm_bridge_write),                    //                                       .write
		.niosii_cpu_spi_mm_bridge_writedata           (niosii_cpu_spi_mm_bridge_writedata),                //                                       .writedata
		.niosii_cpu_spi_mm_bridge_debugaccess         (niosii_cpu_spi_mm_bridge_debugaccess),              //                                       .debugaccess
		.spi_spi_control_port_address                 (mm_interconnect_0_spi_spi_control_port_address),    //                   spi_spi_control_port.address
		.spi_spi_control_port_write                   (mm_interconnect_0_spi_spi_control_port_write),      //                                       .write
		.spi_spi_control_port_read                    (mm_interconnect_0_spi_spi_control_port_read),       //                                       .read
		.spi_spi_control_port_readdata                (mm_interconnect_0_spi_spi_control_port_readdata),   //                                       .readdata
		.spi_spi_control_port_writedata               (mm_interconnect_0_spi_spi_control_port_writedata),  //                                       .writedata
		.spi_spi_control_port_chipselect              (mm_interconnect_0_spi_spi_control_port_chipselect)  //                                       .chipselect
	);

	c5_niosii_spi_slvsec_mm_interconnect_1 mm_interconnect_1 (
		.pll_0_outclk0_clk                                                       (pll_0_outclk0_clk),                                              //                                                     pll_0_outclk0.clk
		.niosii_cpu_reset_reset_bridge_in_reset_reset                            (rst_controller_reset_out_reset),                                 //                            niosii_cpu_reset_reset_bridge_in_reset.reset
		.niosii_cpu_xtrig_mm_bridge_translator_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                 // niosii_cpu_xtrig_mm_bridge_translator_reset_reset_bridge_in_reset.reset
		.niosii_cpu_xtrig_mm_bridge_address                                      (niosii_cpu_xtrig_mm_bridge_address),                             //                                        niosii_cpu_xtrig_mm_bridge.address
		.niosii_cpu_xtrig_mm_bridge_waitrequest                                  (niosii_cpu_xtrig_mm_bridge_waitrequest),                         //                                                                  .waitrequest
		.niosii_cpu_xtrig_mm_bridge_burstcount                                   (niosii_cpu_xtrig_mm_bridge_burstcount),                          //                                                                  .burstcount
		.niosii_cpu_xtrig_mm_bridge_byteenable                                   (niosii_cpu_xtrig_mm_bridge_byteenable),                          //                                                                  .byteenable
		.niosii_cpu_xtrig_mm_bridge_read                                         (niosii_cpu_xtrig_mm_bridge_read),                                //                                                                  .read
		.niosii_cpu_xtrig_mm_bridge_readdata                                     (niosii_cpu_xtrig_mm_bridge_readdata),                            //                                                                  .readdata
		.niosii_cpu_xtrig_mm_bridge_readdatavalid                                (niosii_cpu_xtrig_mm_bridge_readdatavalid),                       //                                                                  .readdatavalid
		.niosii_cpu_xtrig_mm_bridge_write                                        (niosii_cpu_xtrig_mm_bridge_write),                               //                                                                  .write
		.niosii_cpu_xtrig_mm_bridge_writedata                                    (niosii_cpu_xtrig_mm_bridge_writedata),                           //                                                                  .writedata
		.niosii_cpu_xtrig_mm_bridge_debugaccess                                  (niosii_cpu_xtrig_mm_bridge_debugaccess),                         //                                                                  .debugaccess
		.laser_dlp_xtrig_controller_0_avms_address                               (mm_interconnect_1_laser_dlp_xtrig_controller_0_avms_address),    //                                 laser_dlp_xtrig_controller_0_avms.address
		.laser_dlp_xtrig_controller_0_avms_write                                 (mm_interconnect_1_laser_dlp_xtrig_controller_0_avms_write),      //                                                                  .write
		.laser_dlp_xtrig_controller_0_avms_read                                  (mm_interconnect_1_laser_dlp_xtrig_controller_0_avms_read),       //                                                                  .read
		.laser_dlp_xtrig_controller_0_avms_readdata                              (mm_interconnect_1_laser_dlp_xtrig_controller_0_avms_readdata),   //                                                                  .readdata
		.laser_dlp_xtrig_controller_0_avms_writedata                             (mm_interconnect_1_laser_dlp_xtrig_controller_0_avms_writedata),  //                                                                  .writedata
		.laser_dlp_xtrig_controller_0_avms_byteenable                            (mm_interconnect_1_laser_dlp_xtrig_controller_0_avms_byteenable)  //                                                                  .byteenable
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (pll_0_outclk0_clk),              //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
