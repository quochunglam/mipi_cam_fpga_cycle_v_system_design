// c5_niosii_spi_slvsec.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module c5_niosii_spi_slvsec (
		input  wire       clk_clk,                 //        clk.clk
		output wire       inck_en_inck_en_o,       //    inck_en.inck_en_o
		input  wire       key_export,              //        key.export
		output wire [7:0] led_export,              //        led.export
		output wire       reg_1v2_en_reg_1v2_en_o, // reg_1v2_en.reg_1v2_en_o
		output wire       reg_1v8_en_reg_1v8_en_o, // reg_1v8_en.reg_1v8_en_o
		output wire       reg_3v3_en_reg_3v3_en_o, // reg_3v3_en.reg_3v3_en_o
		input  wire       reset_reset_n,           //      reset.reset_n
		input  wire       spi_MISO,                //        spi.MISO
		output wire       spi_MOSI,                //           .MOSI
		output wire       spi_SCLK,                //           .SCLK
		output wire       spi_SS_n,                //           .SS_n
		input  wire [3:0] sw_export,               //         sw.export
		output wire       xclr_xclr_o              //       xclr.xclr_o
	);

	wire         pll_0_outclk0_clk;                                 // pll_0:outclk_0 -> [imx421_poweron:ctrl_clk_i, mm_interconnect_0:pll_0_outclk0_clk, niosii_cpu:clk_clk, rst_controller:clk, spi:clk]
	wire         niosii_cpu_spi_mm_bride_waitrequest;               // mm_interconnect_0:niosii_cpu_spi_mm_bride_waitrequest -> niosii_cpu:spi_mm_bride_waitrequest
	wire  [31:0] niosii_cpu_spi_mm_bride_readdata;                  // mm_interconnect_0:niosii_cpu_spi_mm_bride_readdata -> niosii_cpu:spi_mm_bride_readdata
	wire         niosii_cpu_spi_mm_bride_debugaccess;               // niosii_cpu:spi_mm_bride_debugaccess -> mm_interconnect_0:niosii_cpu_spi_mm_bride_debugaccess
	wire   [9:0] niosii_cpu_spi_mm_bride_address;                   // niosii_cpu:spi_mm_bride_address -> mm_interconnect_0:niosii_cpu_spi_mm_bride_address
	wire         niosii_cpu_spi_mm_bride_read;                      // niosii_cpu:spi_mm_bride_read -> mm_interconnect_0:niosii_cpu_spi_mm_bride_read
	wire   [3:0] niosii_cpu_spi_mm_bride_byteenable;                // niosii_cpu:spi_mm_bride_byteenable -> mm_interconnect_0:niosii_cpu_spi_mm_bride_byteenable
	wire         niosii_cpu_spi_mm_bride_readdatavalid;             // mm_interconnect_0:niosii_cpu_spi_mm_bride_readdatavalid -> niosii_cpu:spi_mm_bride_readdatavalid
	wire  [31:0] niosii_cpu_spi_mm_bride_writedata;                 // niosii_cpu:spi_mm_bride_writedata -> mm_interconnect_0:niosii_cpu_spi_mm_bride_writedata
	wire         niosii_cpu_spi_mm_bride_write;                     // niosii_cpu:spi_mm_bride_write -> mm_interconnect_0:niosii_cpu_spi_mm_bride_write
	wire   [0:0] niosii_cpu_spi_mm_bride_burstcount;                // niosii_cpu:spi_mm_bride_burstcount -> mm_interconnect_0:niosii_cpu_spi_mm_bride_burstcount
	wire         mm_interconnect_0_spi_spi_control_port_chipselect; // mm_interconnect_0:spi_spi_control_port_chipselect -> spi:spi_select
	wire  [15:0] mm_interconnect_0_spi_spi_control_port_readdata;   // spi:data_to_cpu -> mm_interconnect_0:spi_spi_control_port_readdata
	wire   [2:0] mm_interconnect_0_spi_spi_control_port_address;    // mm_interconnect_0:spi_spi_control_port_address -> spi:mem_addr
	wire         mm_interconnect_0_spi_spi_control_port_read;       // mm_interconnect_0:spi_spi_control_port_read -> spi:read_n
	wire         mm_interconnect_0_spi_spi_control_port_write;      // mm_interconnect_0:spi_spi_control_port_write -> spi:write_n
	wire  [15:0] mm_interconnect_0_spi_spi_control_port_writedata;  // mm_interconnect_0:spi_spi_control_port_writedata -> spi:data_from_cpu
	wire         rst_controller_reset_out_reset;                    // rst_controller:reset_out -> [imx421_poweron:ctrl_rst_n_i, mm_interconnect_0:niosii_cpu_reset_reset_bridge_in_reset_reset, mm_interconnect_0:spi_reset_reset_bridge_in_reset_reset, spi:reset_n]

	camera_poweron_sequence_sm #(
		.TIMEOUT_THRESHOLD (34'b0000000000000011110100001001000000)
	) imx421_poweron (
		.ctrl_clk_i   (pll_0_outclk0_clk),               //     clk_in.clk
		.ctrl_rst_n_i (~rst_controller_reset_out_reset), //      rst_n.reset_n
		.reg_1v2_en_o (reg_1v2_en_reg_1v2_en_o),         // reg_1v2_en.reg_1v2_en_o
		.reg_1v8_en_o (reg_1v8_en_reg_1v8_en_o),         // reg_1v8_en.reg_1v8_en_o
		.reg_3v3_en_o (reg_3v3_en_reg_3v3_en_o),         // reg_3v3_en.reg_3v3_en_o
		.inck_en_o    (inck_en_inck_en_o),               //    inck_en.inck_en_o
		.xclr_o       (xclr_xclr_o)                      //       xclr.xclr_o
	);

	c5_niosii_spi_slvsec_niosii_cpu niosii_cpu (
		.clk_clk                    (pll_0_outclk0_clk),                     //          clk.clk
		.key_export                 (key_export),                            //          key.export
		.led_export                 (led_export),                            //          led.export
		.reset_reset_n              (reset_reset_n),                         //        reset.reset_n
		.spi_mm_bride_waitrequest   (niosii_cpu_spi_mm_bride_waitrequest),   // spi_mm_bride.waitrequest
		.spi_mm_bride_readdata      (niosii_cpu_spi_mm_bride_readdata),      //             .readdata
		.spi_mm_bride_readdatavalid (niosii_cpu_spi_mm_bride_readdatavalid), //             .readdatavalid
		.spi_mm_bride_burstcount    (niosii_cpu_spi_mm_bride_burstcount),    //             .burstcount
		.spi_mm_bride_writedata     (niosii_cpu_spi_mm_bride_writedata),     //             .writedata
		.spi_mm_bride_address       (niosii_cpu_spi_mm_bride_address),       //             .address
		.spi_mm_bride_write         (niosii_cpu_spi_mm_bride_write),         //             .write
		.spi_mm_bride_read          (niosii_cpu_spi_mm_bride_read),          //             .read
		.spi_mm_bride_byteenable    (niosii_cpu_spi_mm_bride_byteenable),    //             .byteenable
		.spi_mm_bride_debugaccess   (niosii_cpu_spi_mm_bride_debugaccess),   //             .debugaccess
		.sw_export                  (sw_export)                              //           sw.export
	);

	c5_niosii_spi_slvsec_pll_0 pll_0 (
		.refclk   (clk_clk),           //  refclk.clk
		.rst      (~reset_reset_n),    //   reset.reset
		.outclk_0 (pll_0_outclk0_clk), // outclk0.clk
		.locked   ()                   // (terminated)
	);

	c5_niosii_spi_slvsec_spi spi (
		.clk           (pll_0_outclk0_clk),                                 //              clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                   //            reset.reset_n
		.data_from_cpu (mm_interconnect_0_spi_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_0_spi_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_0_spi_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_0_spi_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_0_spi_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_0_spi_spi_control_port_write),     //                 .write_n
		.irq           (),                                                  //              irq.irq
		.MISO          (spi_MISO),                                          //         external.export
		.MOSI          (spi_MOSI),                                          //                 .export
		.SCLK          (spi_SCLK),                                          //                 .export
		.SS_n          (spi_SS_n)                                           //                 .export
	);

	c5_niosii_spi_slvsec_mm_interconnect_0 mm_interconnect_0 (
		.pll_0_outclk0_clk                            (pll_0_outclk0_clk),                                 //                          pll_0_outclk0.clk
		.niosii_cpu_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                    // niosii_cpu_reset_reset_bridge_in_reset.reset
		.spi_reset_reset_bridge_in_reset_reset        (rst_controller_reset_out_reset),                    //        spi_reset_reset_bridge_in_reset.reset
		.niosii_cpu_spi_mm_bride_address              (niosii_cpu_spi_mm_bride_address),                   //                niosii_cpu_spi_mm_bride.address
		.niosii_cpu_spi_mm_bride_waitrequest          (niosii_cpu_spi_mm_bride_waitrequest),               //                                       .waitrequest
		.niosii_cpu_spi_mm_bride_burstcount           (niosii_cpu_spi_mm_bride_burstcount),                //                                       .burstcount
		.niosii_cpu_spi_mm_bride_byteenable           (niosii_cpu_spi_mm_bride_byteenable),                //                                       .byteenable
		.niosii_cpu_spi_mm_bride_read                 (niosii_cpu_spi_mm_bride_read),                      //                                       .read
		.niosii_cpu_spi_mm_bride_readdata             (niosii_cpu_spi_mm_bride_readdata),                  //                                       .readdata
		.niosii_cpu_spi_mm_bride_readdatavalid        (niosii_cpu_spi_mm_bride_readdatavalid),             //                                       .readdatavalid
		.niosii_cpu_spi_mm_bride_write                (niosii_cpu_spi_mm_bride_write),                     //                                       .write
		.niosii_cpu_spi_mm_bride_writedata            (niosii_cpu_spi_mm_bride_writedata),                 //                                       .writedata
		.niosii_cpu_spi_mm_bride_debugaccess          (niosii_cpu_spi_mm_bride_debugaccess),               //                                       .debugaccess
		.spi_spi_control_port_address                 (mm_interconnect_0_spi_spi_control_port_address),    //                   spi_spi_control_port.address
		.spi_spi_control_port_write                   (mm_interconnect_0_spi_spi_control_port_write),      //                                       .write
		.spi_spi_control_port_read                    (mm_interconnect_0_spi_spi_control_port_read),       //                                       .read
		.spi_spi_control_port_readdata                (mm_interconnect_0_spi_spi_control_port_readdata),   //                                       .readdata
		.spi_spi_control_port_writedata               (mm_interconnect_0_spi_spi_control_port_writedata),  //                                       .writedata
		.spi_spi_control_port_chipselect              (mm_interconnect_0_spi_spi_control_port_chipselect)  //                                       .chipselect
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (pll_0_outclk0_clk),              //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
